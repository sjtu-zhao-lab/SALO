module PE(
  input         clock,
  input         reset,
  input  [8:0]  io_in_q,
  input  [8:0]  io_in_kv,
  input  [4:0]  io_in_inv_sum_exp,
  input  [8:0]  io_in_inv_sum,
  input  [2:0]  io_in_stage,
  output [8:0]  io_out_q,
  output [17:0] io_out_sum,
  output [8:0]  io_out_kv,
  output [2:0]  io_out_stage
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] q; // @[PE.scala 50:16]
  reg [8:0] kv; // @[PE.scala 51:17]
  reg [17:0] sum; // @[PE.scala 52:18]
  reg [2:0] stage; // @[PE.scala 54:20]
  reg [17:0] reg_acc; // @[PE.scala 66:22]
  reg [8:0] reg_prob; // @[PE.scala 67:23]
  reg [4:0] reg_max_exp; // @[PE.scala 75:26]
  wire [4:0] integer_bits = reg_acc[15:11]; // @[PE.scala 88:43]
  wire [8:0] fraction_bits = {1'b0,$signed(reg_acc[10:3])}; // @[PE.scala 89:41]
  wire [8:0] _GEN_1 = 2'h1 == fraction_bits[7:6] ? $signed(9'she) : $signed(9'shc); // @[PE.scala 90:7 PE.scala 90:7]
  wire [8:0] _GEN_2 = 2'h2 == fraction_bits[7:6] ? $signed(9'sh11) : $signed(_GEN_1); // @[PE.scala 90:7 PE.scala 90:7]
  wire [8:0] k = 2'h3 == fraction_bits[7:6] ? $signed(9'sh14) : $signed(_GEN_2); // @[PE.scala 90:7 PE.scala 90:7]
  wire [17:0] _GEN_5 = 2'h1 == fraction_bits[7:6] ? $signed(18'shf6) : $signed(18'shff); // @[PE.scala 91:7 PE.scala 91:7]
  wire [17:0] _GEN_6 = 2'h2 == fraction_bits[7:6] ? $signed(18'she1) : $signed(_GEN_5); // @[PE.scala 91:7 PE.scala 91:7]
  wire [17:0] b = 2'h3 == fraction_bits[7:6] ? $signed(18'shb9) : $signed(_GEN_6); // @[PE.scala 91:7 PE.scala 91:7]
  wire  _T_2 = ~reset; // @[PE.scala 92:11]
  wire [8:0] _T_4 = {1'b0,$signed(reg_acc[8:1])}; // @[PE.scala 103:51]
  wire [8:0] _oprand1_T_4 = 3'h0 == io_in_stage ? $signed(io_in_q) : $signed(9'sh0); // @[Mux.scala 80:57]
  wire [8:0] _oprand1_T_6 = 3'h1 == io_in_stage ? $signed(k) : $signed(_oprand1_T_4); // @[Mux.scala 80:57]
  wire [8:0] _oprand1_T_8 = 3'h3 == io_in_stage ? $signed(_T_4) : $signed(_oprand1_T_6); // @[Mux.scala 80:57]
  wire [8:0] oprand1 = 3'h4 == io_in_stage ? $signed(reg_prob) : $signed(_oprand1_T_8); // @[Mux.scala 80:57]
  wire [8:0] _oprand2_T_2 = 3'h0 == io_in_stage ? $signed(io_in_kv) : $signed(9'sh0); // @[Mux.scala 80:57]
  wire [8:0] _oprand2_T_4 = 3'h1 == io_in_stage ? $signed(fraction_bits) : $signed(_oprand2_T_2); // @[Mux.scala 80:57]
  wire [8:0] _oprand2_T_6 = 3'h3 == io_in_stage ? $signed(io_in_inv_sum) : $signed(_oprand2_T_4); // @[Mux.scala 80:57]
  wire [8:0] oprand2 = 3'h4 == io_in_stage ? $signed(io_in_kv) : $signed(_oprand2_T_6); // @[Mux.scala 80:57]
  wire [17:0] _oprand3_T_1 = 3'h0 == io_in_stage ? $signed(reg_acc) : $signed(18'sh0); // @[Mux.scala 80:57]
  wire [17:0] _oprand3_T_3 = 3'h1 == io_in_stage ? $signed(b) : $signed(_oprand3_T_1); // @[Mux.scala 80:57]
  wire [17:0] _oprand3_T_5 = 3'h2 == io_in_stage ? $signed(18'sh0) : $signed(_oprand3_T_3); // @[Mux.scala 80:57]
  wire [17:0] _oprand3_T_7 = 3'h3 == io_in_stage ? $signed(18'sh0) : $signed(_oprand3_T_5); // @[Mux.scala 80:57]
  wire [17:0] oprand3 = 3'h4 == io_in_stage ? $signed(18'sh0) : $signed(_oprand3_T_7); // @[Mux.scala 80:57]
  wire  _product_T = io_in_stage == 3'h2; // @[PE.scala 111:31]
  wire [17:0] _product_T_1 = $signed(oprand1) * $signed(oprand2); // @[PE.scala 111:60]
  wire [17:0] product = io_in_stage == 3'h2 ? $signed(18'sh0) : $signed(_product_T_1); // @[PE.scala 111:19]
  wire  _oprand4_T = io_in_stage == 3'h4; // @[PE.scala 112:31]
  wire [14:0] _oprand4_T_1 = product[17:3]; // @[PE.scala 112:47]
  wire  _oprand4_T_2 = io_in_stage == 3'h1; // @[PE.scala 112:68]
  wire [13:0] _oprand4_T_3 = product[17:4]; // @[PE.scala 112:84]
  wire [17:0] _oprand4_T_4 = io_in_stage == 3'h1 ? $signed({{4{_oprand4_T_3[13]}},_oprand4_T_3}) : $signed(product); // @[PE.scala 112:56]
  wire [17:0] oprand4 = io_in_stage == 3'h4 ? $signed({{3{_oprand4_T_1[14]}},_oprand4_T_1}) : $signed(_oprand4_T_4); // @[PE.scala 112:19]
  wire [17:0] result = $signed(oprand3) + $signed(oprand4); // @[PE.scala 113:23]
  wire [4:0] _reg_prob_T_3 = $signed(io_in_inv_sum_exp) - $signed(reg_max_exp); // @[PE.scala 150:72]
  wire [17:0] _reg_prob_T_4 = $signed(result) >>> _reg_prob_T_3; // @[PE.scala 150:29]
  wire [8:0] _reg_prob_T_6 = _reg_prob_T_4[15:7]; // @[PE.scala 150:94]
  assign io_out_q = q; // @[PE.scala 60:14]
  assign io_out_sum = sum; // @[PE.scala 62:16]
  assign io_out_kv = kv; // @[PE.scala 61:15]
  assign io_out_stage = stage; // @[PE.scala 64:18]
  always @(posedge clock) begin
    q <= io_in_q; // @[PE.scala 56:7]
    kv <= io_in_kv; // @[PE.scala 57:8]
    if (_product_T) begin // @[PE.scala 131:35]
      sum <= result; // @[PE.scala 146:13]
    end else if (_oprand4_T) begin // @[PE.scala 154:35]
      sum <= result; // @[PE.scala 158:13]
    end
    stage <= io_in_stage; // @[PE.scala 58:11]
    if (io_in_stage == 3'h0) begin // @[PE.scala 119:29]
      reg_acc <= result; // @[PE.scala 120:17]
    end else if (_oprand4_T_2) begin // @[PE.scala 125:35]
      reg_acc <= result; // @[PE.scala 126:17]
    end else if (_product_T) begin // @[PE.scala 131:35]
      reg_acc <= 18'sh0; // @[PE.scala 143:17]
    end
    if (io_in_stage == 3'h3) begin // @[PE.scala 148:35]
      reg_prob <= _reg_prob_T_6; // @[PE.scala 150:18]
    end
    if (_oprand4_T_2) begin // @[PE.scala 125:35]
      reg_max_exp <= integer_bits; // @[PE.scala 128:21]
    end else if (_product_T) begin // @[PE.scala 131:35]
      reg_max_exp <= 5'sh0; // @[PE.scala 145:21]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"reg_acc = %b\n",reg_acc); // @[PE.scala 92:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2) begin
          $fwrite(32'h80000002,"ext_acc = %b\n",{1'b0,$signed(reg_acc[8:1])}); // @[PE.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2) begin
          $fwrite(32'h80000002,"inv_sum = %b\n",io_in_inv_sum); // @[PE.scala 104:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2) begin
          $fwrite(32'h80000002,"reg_prob = %b\n",reg_prob); // @[PE.scala 105:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  q = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  kv = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  sum = _RAND_2[17:0];
  _RAND_3 = {1{`RANDOM}};
  stage = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  reg_acc = _RAND_4[17:0];
  _RAND_5 = {1{`RANDOM}};
  reg_prob = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  reg_max_exp = _RAND_6[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PE_1(
  input         clock,
  input         reset,
  input  [8:0]  io_in_q,
  input  [17:0] io_in_sum,
  input  [4:0]  io_in_sum_exp,
  input  [8:0]  io_in_kv,
  input  [4:0]  io_in_inv_sum_exp,
  input  [8:0]  io_in_inv_sum,
  input  [2:0]  io_in_stage,
  output [8:0]  io_out_q,
  output [17:0] io_out_sum,
  output [4:0]  io_out_sum_exp,
  output [8:0]  io_out_kv,
  output [2:0]  io_out_stage
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] q; // @[PE.scala 50:16]
  reg [8:0] kv; // @[PE.scala 51:17]
  reg [17:0] sum; // @[PE.scala 52:18]
  reg [4:0] sum_exp; // @[PE.scala 53:22]
  reg [2:0] stage; // @[PE.scala 54:20]
  reg [17:0] reg_acc; // @[PE.scala 66:22]
  reg [8:0] reg_prob; // @[PE.scala 67:23]
  reg [4:0] reg_max_exp; // @[PE.scala 75:26]
  wire [4:0] integer_bits = reg_acc[15:11]; // @[PE.scala 88:43]
  wire [8:0] fraction_bits = {1'b0,$signed(reg_acc[10:3])}; // @[PE.scala 89:41]
  wire [8:0] _GEN_1 = 2'h1 == fraction_bits[7:6] ? $signed(9'she) : $signed(9'shc); // @[PE.scala 90:7 PE.scala 90:7]
  wire [8:0] _GEN_2 = 2'h2 == fraction_bits[7:6] ? $signed(9'sh11) : $signed(_GEN_1); // @[PE.scala 90:7 PE.scala 90:7]
  wire [8:0] k = 2'h3 == fraction_bits[7:6] ? $signed(9'sh14) : $signed(_GEN_2); // @[PE.scala 90:7 PE.scala 90:7]
  wire [17:0] _GEN_5 = 2'h1 == fraction_bits[7:6] ? $signed(18'shf6) : $signed(18'shff); // @[PE.scala 91:7 PE.scala 91:7]
  wire [17:0] _GEN_6 = 2'h2 == fraction_bits[7:6] ? $signed(18'she1) : $signed(_GEN_5); // @[PE.scala 91:7 PE.scala 91:7]
  wire [17:0] b = 2'h3 == fraction_bits[7:6] ? $signed(18'shb9) : $signed(_GEN_6); // @[PE.scala 91:7 PE.scala 91:7]
  wire  _T_2 = ~reset; // @[PE.scala 92:11]
  wire [8:0] _T_4 = {1'b0,$signed(reg_acc[8:1])}; // @[PE.scala 103:51]
  wire [8:0] _oprand1_T_4 = 3'h0 == io_in_stage ? $signed(io_in_q) : $signed(9'sh0); // @[Mux.scala 80:57]
  wire [8:0] _oprand1_T_6 = 3'h1 == io_in_stage ? $signed(k) : $signed(_oprand1_T_4); // @[Mux.scala 80:57]
  wire [8:0] _oprand1_T_8 = 3'h3 == io_in_stage ? $signed(_T_4) : $signed(_oprand1_T_6); // @[Mux.scala 80:57]
  wire [8:0] oprand1 = 3'h4 == io_in_stage ? $signed(reg_prob) : $signed(_oprand1_T_8); // @[Mux.scala 80:57]
  wire [8:0] _oprand2_T_2 = 3'h0 == io_in_stage ? $signed(io_in_kv) : $signed(9'sh0); // @[Mux.scala 80:57]
  wire [8:0] _oprand2_T_4 = 3'h1 == io_in_stage ? $signed(fraction_bits) : $signed(_oprand2_T_2); // @[Mux.scala 80:57]
  wire [8:0] _oprand2_T_6 = 3'h3 == io_in_stage ? $signed(io_in_inv_sum) : $signed(_oprand2_T_4); // @[Mux.scala 80:57]
  wire [8:0] oprand2 = 3'h4 == io_in_stage ? $signed(io_in_kv) : $signed(_oprand2_T_6); // @[Mux.scala 80:57]
  wire [17:0] _oprand3_T_1 = 3'h0 == io_in_stage ? $signed(reg_acc) : $signed(18'sh0); // @[Mux.scala 80:57]
  wire [17:0] _oprand3_T_3 = 3'h1 == io_in_stage ? $signed(b) : $signed(_oprand3_T_1); // @[Mux.scala 80:57]
  wire  _T_14 = io_in_stage == 3'h1; // @[PE.scala 125:27]
  wire  _T_15 = io_in_stage == 3'h2; // @[PE.scala 131:27]
  wire [4:0] _shifted_sum_T_3 = $signed(reg_max_exp) - $signed(io_in_sum_exp); // @[PE.scala 139:81]
  wire [17:0] _shifted_sum_T_4 = $signed(io_in_sum) >>> _shifted_sum_T_3; // @[PE.scala 139:42]
  wire [17:0] shifted_sum = $signed(reg_max_exp) < $signed(io_in_sum_exp) ? $signed(io_in_sum) : $signed(
    _shifted_sum_T_4); // @[PE.scala 133:47 PE.scala 135:29 PE.scala 139:29]
  wire [17:0] _oprand3_T_5 = 3'h2 == io_in_stage ? $signed(shifted_sum) : $signed(_oprand3_T_3); // @[Mux.scala 80:57]
  wire [17:0] _oprand3_T_7 = 3'h3 == io_in_stage ? $signed(18'sh0) : $signed(_oprand3_T_5); // @[Mux.scala 80:57]
  wire [17:0] oprand3 = 3'h4 == io_in_stage ? $signed(io_in_sum) : $signed(_oprand3_T_7); // @[Mux.scala 80:57]
  wire [17:0] _product_T_1 = $signed(oprand1) * $signed(oprand2); // @[PE.scala 111:60]
  wire [4:0] _shifted_acc_T_3 = $signed(io_in_sum_exp) - $signed(reg_max_exp); // @[PE.scala 134:79]
  wire [17:0] _shifted_acc_T_4 = $signed(reg_acc) >>> _shifted_acc_T_3; // @[PE.scala 134:40]
  wire [17:0] shifted_acc = $signed(reg_max_exp) < $signed(io_in_sum_exp) ? $signed(_shifted_acc_T_4) : $signed(reg_acc)
    ; // @[PE.scala 133:47 PE.scala 134:29 PE.scala 138:29]
  wire [17:0] product = _T_15 ? $signed(shifted_acc) : $signed(_product_T_1); // @[PE.scala 111:19]
  wire  _oprand4_T = io_in_stage == 3'h4; // @[PE.scala 112:31]
  wire [14:0] _oprand4_T_1 = product[17:3]; // @[PE.scala 112:47]
  wire [13:0] _oprand4_T_3 = product[17:4]; // @[PE.scala 112:84]
  wire [17:0] _oprand4_T_4 = _T_14 ? $signed({{4{_oprand4_T_3[13]}},_oprand4_T_3}) : $signed(product); // @[PE.scala 112:56]
  wire [17:0] oprand4 = io_in_stage == 3'h4 ? $signed({{3{_oprand4_T_1[14]}},_oprand4_T_1}) : $signed(_oprand4_T_4); // @[PE.scala 112:19]
  wire [17:0] result = $signed(oprand3) + $signed(oprand4); // @[PE.scala 113:23]
  wire [4:0] _reg_prob_T_3 = $signed(io_in_inv_sum_exp) - $signed(reg_max_exp); // @[PE.scala 150:72]
  wire [17:0] _reg_prob_T_4 = $signed(result) >>> _reg_prob_T_3; // @[PE.scala 150:29]
  wire [8:0] _reg_prob_T_6 = _reg_prob_T_4[15:7]; // @[PE.scala 150:94]
  assign io_out_q = q; // @[PE.scala 60:14]
  assign io_out_sum = sum; // @[PE.scala 62:16]
  assign io_out_sum_exp = sum_exp; // @[PE.scala 63:20]
  assign io_out_kv = kv; // @[PE.scala 61:15]
  assign io_out_stage = stage; // @[PE.scala 64:18]
  always @(posedge clock) begin
    q <= io_in_q; // @[PE.scala 56:7]
    kv <= io_in_kv; // @[PE.scala 57:8]
    if (io_in_stage == 3'h2) begin // @[PE.scala 131:35]
      sum <= result; // @[PE.scala 146:13]
    end else if (_oprand4_T) begin // @[PE.scala 154:35]
      sum <= result; // @[PE.scala 158:13]
    end
    if (io_in_stage == 3'h2) begin // @[PE.scala 131:35]
      if ($signed(reg_max_exp) < $signed(io_in_sum_exp)) begin // @[PE.scala 133:47]
        sum_exp <= io_in_sum_exp; // @[PE.scala 136:25]
      end else begin
        sum_exp <= reg_max_exp; // @[PE.scala 140:25]
      end
    end
    stage <= io_in_stage; // @[PE.scala 58:11]
    if (io_in_stage == 3'h0) begin // @[PE.scala 119:29]
      reg_acc <= result; // @[PE.scala 120:17]
    end else if (io_in_stage == 3'h1) begin // @[PE.scala 125:35]
      reg_acc <= result; // @[PE.scala 126:17]
    end else if (io_in_stage == 3'h2) begin // @[PE.scala 131:35]
      if ($signed(reg_max_exp) < $signed(io_in_sum_exp)) begin // @[PE.scala 133:47]
        reg_acc <= _shifted_acc_T_4; // @[PE.scala 134:29]
      end
    end
    if (io_in_stage == 3'h3) begin // @[PE.scala 148:35]
      reg_prob <= _reg_prob_T_6; // @[PE.scala 150:18]
    end
    if (io_in_stage == 3'h1) begin // @[PE.scala 125:35]
      reg_max_exp <= integer_bits; // @[PE.scala 128:21]
    end else if (io_in_stage == 3'h2) begin // @[PE.scala 131:35]
      if ($signed(reg_max_exp) < $signed(io_in_sum_exp)) begin // @[PE.scala 133:47]
        reg_max_exp <= io_in_sum_exp; // @[PE.scala 136:25]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset) begin
          $fwrite(32'h80000002,"reg_acc = %b\n",reg_acc); // @[PE.scala 92:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2) begin
          $fwrite(32'h80000002,"ext_acc = %b\n",{1'b0,$signed(reg_acc[8:1])}); // @[PE.scala 103:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2) begin
          $fwrite(32'h80000002,"inv_sum = %b\n",io_in_inv_sum); // @[PE.scala 104:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2) begin
          $fwrite(32'h80000002,"reg_prob = %b\n",reg_prob); // @[PE.scala 105:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  q = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  kv = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  sum = _RAND_2[17:0];
  _RAND_3 = {1{`RANDOM}};
  sum_exp = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  stage = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  reg_acc = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  reg_prob = _RAND_6[8:0];
  _RAND_7 = {1{`RANDOM}};
  reg_max_exp = _RAND_7[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module InverseModule(
  input  [17:0] io_in_sum,
  input  [4:0]  io_in_exp,
  output [8:0]  io_out_inv_sum,
  output [4:0]  io_out_inv_sum_exp
);
  wire [17:0] _io_out_inv_sum_T_1 = 18'h20000 / io_in_sum; // @[InverseModule.scala 20:35]
  wire [8:0] _io_out_inv_sum_T_3 = _io_out_inv_sum_T_1[17:9]; // @[InverseModule.scala 20:75]
  wire [4:0] _GEN_0 = _io_out_inv_sum_T_3[8:4]; // @[InverseModule.scala 20:20]
  assign io_out_inv_sum = {{4{_GEN_0[4]}},_GEN_0}; // @[InverseModule.scala 20:20]
  assign io_out_inv_sum_exp = io_in_exp; // @[InverseModule.scala 21:24]
endmodule
module WeightedSumModule(
  input         clock,
  input         reset,
  input  [17:0] io_in_sum,
  input  [4:0]  io_in_exp,
  input  [1:0]  io_control,
  output [17:0] io_out_port
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
`endif // RANDOMIZE_REG_INIT
  reg [17:0] sum; // @[WeightedSumModule.scala 21:18]
  reg [4:0] exp; // @[WeightedSumModule.scala 22:18]
  reg [17:0] c; // @[WeightedSumModule.scala 23:17]
  reg [4:0] c_exp; // @[WeightedSumModule.scala 24:20]
  reg [17:0] w1; // @[WeightedSumModule.scala 26:17]
  reg [17:0] w2; // @[WeightedSumModule.scala 27:17]
  reg [17:0] buffer_0; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_1; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_2; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_3; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_4; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_5; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_6; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_7; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_8; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_9; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_10; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_11; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_12; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_13; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_14; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_15; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_16; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_17; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_18; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_19; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_20; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_21; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_22; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_23; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_24; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_25; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_26; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_27; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_28; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_29; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_30; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_31; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_32; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_33; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_34; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_35; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_36; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_37; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_38; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_39; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_40; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_41; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_42; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_43; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_44; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_45; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_46; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_47; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_48; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_49; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_50; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_51; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_52; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_53; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_54; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_55; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_56; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_57; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_58; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_59; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_60; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_61; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_62; // @[WeightedSumModule.scala 28:21]
  reg [17:0] buffer_63; // @[WeightedSumModule.scala 28:21]
  wire  _T = io_control == 2'h3; // @[WeightedSumModule.scala 29:42]
  reg [5:0] cnt; // @[Counter.scala 60:40]
  wire [5:0] _wrap_value_T_1 = cnt + 6'h1; // @[Counter.scala 76:24]
  wire [4:0] _shifted_sum_T_3 = $signed(io_in_exp) - $signed(exp); // @[WeightedSumModule.scala 48:59]
  wire [17:0] _shifted_sum_T_4 = $signed(sum) >>> _shifted_sum_T_3; // @[WeightedSumModule.scala 48:32]
  wire [4:0] _shifted_in_sum_T_3 = $signed(exp) - $signed(io_in_exp); // @[WeightedSumModule.scala 53:68]
  wire [17:0] _shifted_in_sum_T_4 = $signed(io_in_sum) >>> _shifted_in_sum_T_3; // @[WeightedSumModule.scala 53:41]
  wire [17:0] shifted_sum = $signed(exp) < $signed(io_in_exp) ? $signed(_shifted_sum_T_4) : $signed(sum); // @[WeightedSumModule.scala 47:31 WeightedSumModule.scala 48:25 WeightedSumModule.scala 52:25]
  wire [17:0] shifted_in_sum = $signed(exp) < $signed(io_in_exp) ? $signed(io_in_sum) : $signed(_shifted_in_sum_T_4); // @[WeightedSumModule.scala 47:31 WeightedSumModule.scala 49:28 WeightedSumModule.scala 53:28]
  wire [17:0] _c_T_2 = $signed(shifted_sum) + $signed(shifted_in_sum); // @[WeightedSumModule.scala 56:26]
  wire [21:0] _w1_T_1 = {$signed(w1), 4'h0}; // @[WeightedSumModule.scala 64:33]
  wire [21:0] _w1_T_3 = _w1_T_1 / c; // @[WeightedSumModule.scala 64:36]
  wire [17:0] _w1_T_5 = _w1_T_3[21:4]; // @[WeightedSumModule.scala 64:68]
  wire [21:0] _w2_T_1 = {$signed(w2), 4'h0}; // @[WeightedSumModule.scala 65:33]
  wire [21:0] _w2_T_3 = _w2_T_1 / c; // @[WeightedSumModule.scala 65:36]
  wire [17:0] _w2_T_5 = _w2_T_3[21:4]; // @[WeightedSumModule.scala 65:68]
  wire [17:0] _GEN_6 = 6'h1 == cnt ? $signed(buffer_1) : $signed(buffer_0); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_7 = 6'h2 == cnt ? $signed(buffer_2) : $signed(_GEN_6); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_8 = 6'h3 == cnt ? $signed(buffer_3) : $signed(_GEN_7); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_9 = 6'h4 == cnt ? $signed(buffer_4) : $signed(_GEN_8); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_10 = 6'h5 == cnt ? $signed(buffer_5) : $signed(_GEN_9); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_11 = 6'h6 == cnt ? $signed(buffer_6) : $signed(_GEN_10); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_12 = 6'h7 == cnt ? $signed(buffer_7) : $signed(_GEN_11); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_13 = 6'h8 == cnt ? $signed(buffer_8) : $signed(_GEN_12); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_14 = 6'h9 == cnt ? $signed(buffer_9) : $signed(_GEN_13); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_15 = 6'ha == cnt ? $signed(buffer_10) : $signed(_GEN_14); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_16 = 6'hb == cnt ? $signed(buffer_11) : $signed(_GEN_15); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_17 = 6'hc == cnt ? $signed(buffer_12) : $signed(_GEN_16); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_18 = 6'hd == cnt ? $signed(buffer_13) : $signed(_GEN_17); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_19 = 6'he == cnt ? $signed(buffer_14) : $signed(_GEN_18); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_20 = 6'hf == cnt ? $signed(buffer_15) : $signed(_GEN_19); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_21 = 6'h10 == cnt ? $signed(buffer_16) : $signed(_GEN_20); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_22 = 6'h11 == cnt ? $signed(buffer_17) : $signed(_GEN_21); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_23 = 6'h12 == cnt ? $signed(buffer_18) : $signed(_GEN_22); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_24 = 6'h13 == cnt ? $signed(buffer_19) : $signed(_GEN_23); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_25 = 6'h14 == cnt ? $signed(buffer_20) : $signed(_GEN_24); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_26 = 6'h15 == cnt ? $signed(buffer_21) : $signed(_GEN_25); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_27 = 6'h16 == cnt ? $signed(buffer_22) : $signed(_GEN_26); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_28 = 6'h17 == cnt ? $signed(buffer_23) : $signed(_GEN_27); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_29 = 6'h18 == cnt ? $signed(buffer_24) : $signed(_GEN_28); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_30 = 6'h19 == cnt ? $signed(buffer_25) : $signed(_GEN_29); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_31 = 6'h1a == cnt ? $signed(buffer_26) : $signed(_GEN_30); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_32 = 6'h1b == cnt ? $signed(buffer_27) : $signed(_GEN_31); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_33 = 6'h1c == cnt ? $signed(buffer_28) : $signed(_GEN_32); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_34 = 6'h1d == cnt ? $signed(buffer_29) : $signed(_GEN_33); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_35 = 6'h1e == cnt ? $signed(buffer_30) : $signed(_GEN_34); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_36 = 6'h1f == cnt ? $signed(buffer_31) : $signed(_GEN_35); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_37 = 6'h20 == cnt ? $signed(buffer_32) : $signed(_GEN_36); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_38 = 6'h21 == cnt ? $signed(buffer_33) : $signed(_GEN_37); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_39 = 6'h22 == cnt ? $signed(buffer_34) : $signed(_GEN_38); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_40 = 6'h23 == cnt ? $signed(buffer_35) : $signed(_GEN_39); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_41 = 6'h24 == cnt ? $signed(buffer_36) : $signed(_GEN_40); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_42 = 6'h25 == cnt ? $signed(buffer_37) : $signed(_GEN_41); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_43 = 6'h26 == cnt ? $signed(buffer_38) : $signed(_GEN_42); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_44 = 6'h27 == cnt ? $signed(buffer_39) : $signed(_GEN_43); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_45 = 6'h28 == cnt ? $signed(buffer_40) : $signed(_GEN_44); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_46 = 6'h29 == cnt ? $signed(buffer_41) : $signed(_GEN_45); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_47 = 6'h2a == cnt ? $signed(buffer_42) : $signed(_GEN_46); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_48 = 6'h2b == cnt ? $signed(buffer_43) : $signed(_GEN_47); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_49 = 6'h2c == cnt ? $signed(buffer_44) : $signed(_GEN_48); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_50 = 6'h2d == cnt ? $signed(buffer_45) : $signed(_GEN_49); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_51 = 6'h2e == cnt ? $signed(buffer_46) : $signed(_GEN_50); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_52 = 6'h2f == cnt ? $signed(buffer_47) : $signed(_GEN_51); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_53 = 6'h30 == cnt ? $signed(buffer_48) : $signed(_GEN_52); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_54 = 6'h31 == cnt ? $signed(buffer_49) : $signed(_GEN_53); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_55 = 6'h32 == cnt ? $signed(buffer_50) : $signed(_GEN_54); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_56 = 6'h33 == cnt ? $signed(buffer_51) : $signed(_GEN_55); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_57 = 6'h34 == cnt ? $signed(buffer_52) : $signed(_GEN_56); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_58 = 6'h35 == cnt ? $signed(buffer_53) : $signed(_GEN_57); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_59 = 6'h36 == cnt ? $signed(buffer_54) : $signed(_GEN_58); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_60 = 6'h37 == cnt ? $signed(buffer_55) : $signed(_GEN_59); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_61 = 6'h38 == cnt ? $signed(buffer_56) : $signed(_GEN_60); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_62 = 6'h39 == cnt ? $signed(buffer_57) : $signed(_GEN_61); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_63 = 6'h3a == cnt ? $signed(buffer_58) : $signed(_GEN_62); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_64 = 6'h3b == cnt ? $signed(buffer_59) : $signed(_GEN_63); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_65 = 6'h3c == cnt ? $signed(buffer_60) : $signed(_GEN_64); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_66 = 6'h3d == cnt ? $signed(buffer_61) : $signed(_GEN_65); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_67 = 6'h3e == cnt ? $signed(buffer_62) : $signed(_GEN_66); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [17:0] _GEN_68 = 6'h3f == cnt ? $signed(buffer_63) : $signed(_GEN_67); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  wire [35:0] _buffer_T = $signed(w1) * $signed(_GEN_68); // @[WeightedSumModule.scala 72:27]
  wire [35:0] _buffer_T_1 = $signed(w2) * $signed(io_in_sum); // @[WeightedSumModule.scala 72:46]
  wire [35:0] _buffer_T_4 = $signed(_buffer_T) + $signed(_buffer_T_1); // @[WeightedSumModule.scala 72:41]
  wire [27:0] _GEN_415 = _buffer_T_4[35:8]; // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21]
  wire [17:0] _buffer_cnt_0 = _GEN_415[17:0]; // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21]
  wire [17:0] _GEN_69 = 6'h0 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_0); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_70 = 6'h1 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_1); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_71 = 6'h2 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_2); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_72 = 6'h3 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_3); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_73 = 6'h4 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_4); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_74 = 6'h5 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_5); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_75 = 6'h6 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_6); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_76 = 6'h7 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_7); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_77 = 6'h8 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_8); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_78 = 6'h9 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_9); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_79 = 6'ha == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_10); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_80 = 6'hb == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_11); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_81 = 6'hc == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_12); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_82 = 6'hd == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_13); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_83 = 6'he == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_14); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_84 = 6'hf == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_15); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_85 = 6'h10 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_16); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_86 = 6'h11 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_17); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_87 = 6'h12 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_18); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_88 = 6'h13 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_19); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_89 = 6'h14 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_20); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_90 = 6'h15 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_21); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_91 = 6'h16 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_22); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_92 = 6'h17 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_23); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_93 = 6'h18 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_24); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_94 = 6'h19 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_25); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_95 = 6'h1a == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_26); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_96 = 6'h1b == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_27); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_97 = 6'h1c == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_28); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_98 = 6'h1d == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_29); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_99 = 6'h1e == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_30); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_100 = 6'h1f == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_31); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_101 = 6'h20 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_32); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_102 = 6'h21 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_33); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_103 = 6'h22 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_34); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_104 = 6'h23 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_35); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_105 = 6'h24 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_36); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_106 = 6'h25 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_37); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_107 = 6'h26 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_38); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_108 = 6'h27 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_39); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_109 = 6'h28 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_40); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_110 = 6'h29 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_41); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_111 = 6'h2a == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_42); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_112 = 6'h2b == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_43); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_113 = 6'h2c == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_44); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_114 = 6'h2d == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_45); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_115 = 6'h2e == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_46); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_116 = 6'h2f == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_47); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_117 = 6'h30 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_48); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_118 = 6'h31 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_49); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_119 = 6'h32 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_50); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_120 = 6'h33 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_51); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_121 = 6'h34 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_52); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_122 = 6'h35 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_53); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_123 = 6'h36 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_54); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_124 = 6'h37 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_55); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_125 = 6'h38 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_56); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_126 = 6'h39 == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_57); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_127 = 6'h3a == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_58); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_128 = 6'h3b == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_59); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_129 = 6'h3c == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_60); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_130 = 6'h3d == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_61); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_131 = 6'h3e == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_62); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  wire [17:0] _GEN_132 = 6'h3f == cnt ? $signed(_buffer_cnt_0) : $signed(buffer_63); // @[WeightedSumModule.scala 72:21 WeightedSumModule.scala 72:21 WeightedSumModule.scala 28:21]
  assign io_out_port = 6'h3f == cnt ? $signed(buffer_63) : $signed(_GEN_67); // @[WeightedSumModule.scala 72:27 WeightedSumModule.scala 72:27]
  always @(posedge clock) begin
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      sum <= 18'sh0; // @[WeightedSumModule.scala 44:13]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (io_control == 2'h2) begin // @[WeightedSumModule.scala 63:33]
        sum <= c; // @[WeightedSumModule.scala 66:13]
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      exp <= 5'sh0; // @[WeightedSumModule.scala 45:13]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (io_control == 2'h2) begin // @[WeightedSumModule.scala 63:33]
        exp <= c_exp; // @[WeightedSumModule.scala 67:13]
      end
    end
    if (!(io_control == 2'h0)) begin // @[WeightedSumModule.scala 40:27]
      if (io_control == 2'h1) begin // @[WeightedSumModule.scala 46:33]
        c <= _c_T_2; // @[WeightedSumModule.scala 56:11]
      end
    end
    if (!(io_control == 2'h0)) begin // @[WeightedSumModule.scala 40:27]
      if (io_control == 2'h1) begin // @[WeightedSumModule.scala 46:33]
        if ($signed(exp) < $signed(io_in_exp)) begin // @[WeightedSumModule.scala 47:31]
          c_exp <= io_in_exp; // @[WeightedSumModule.scala 50:21]
        end else begin
          c_exp <= exp; // @[WeightedSumModule.scala 54:21]
        end
      end
    end
    if (!(io_control == 2'h0)) begin // @[WeightedSumModule.scala 40:27]
      if (io_control == 2'h1) begin // @[WeightedSumModule.scala 46:33]
        if ($signed(exp) < $signed(io_in_exp)) begin // @[WeightedSumModule.scala 47:31]
          w1 <= _shifted_sum_T_4; // @[WeightedSumModule.scala 48:25]
        end else begin
          w1 <= sum; // @[WeightedSumModule.scala 52:25]
        end
      end else if (io_control == 2'h2) begin // @[WeightedSumModule.scala 63:33]
        w1 <= _w1_T_5; // @[WeightedSumModule.scala 64:12]
      end
    end
    if (!(io_control == 2'h0)) begin // @[WeightedSumModule.scala 40:27]
      if (io_control == 2'h1) begin // @[WeightedSumModule.scala 46:33]
        if ($signed(exp) < $signed(io_in_exp)) begin // @[WeightedSumModule.scala 47:31]
          w2 <= io_in_sum; // @[WeightedSumModule.scala 49:28]
        end else begin
          w2 <= _shifted_in_sum_T_4; // @[WeightedSumModule.scala 53:28]
        end
      end else if (io_control == 2'h2) begin // @[WeightedSumModule.scala 63:33]
        w2 <= _w2_T_5; // @[WeightedSumModule.scala 65:12]
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_0 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_0 <= _GEN_69;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_1 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_1 <= _GEN_70;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_2 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_2 <= _GEN_71;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_3 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_3 <= _GEN_72;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_4 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_4 <= _GEN_73;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_5 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_5 <= _GEN_74;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_6 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_6 <= _GEN_75;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_7 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_7 <= _GEN_76;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_8 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_8 <= _GEN_77;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_9 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_9 <= _GEN_78;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_10 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_10 <= _GEN_79;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_11 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_11 <= _GEN_80;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_12 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_12 <= _GEN_81;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_13 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_13 <= _GEN_82;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_14 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_14 <= _GEN_83;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_15 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_15 <= _GEN_84;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_16 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_16 <= _GEN_85;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_17 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_17 <= _GEN_86;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_18 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_18 <= _GEN_87;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_19 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_19 <= _GEN_88;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_20 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_20 <= _GEN_89;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_21 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_21 <= _GEN_90;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_22 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_22 <= _GEN_91;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_23 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_23 <= _GEN_92;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_24 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_24 <= _GEN_93;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_25 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_25 <= _GEN_94;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_26 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_26 <= _GEN_95;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_27 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_27 <= _GEN_96;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_28 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_28 <= _GEN_97;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_29 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_29 <= _GEN_98;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_30 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_30 <= _GEN_99;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_31 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_31 <= _GEN_100;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_32 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_32 <= _GEN_101;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_33 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_33 <= _GEN_102;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_34 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_34 <= _GEN_103;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_35 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_35 <= _GEN_104;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_36 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_36 <= _GEN_105;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_37 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_37 <= _GEN_106;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_38 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_38 <= _GEN_107;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_39 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_39 <= _GEN_108;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_40 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_40 <= _GEN_109;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_41 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_41 <= _GEN_110;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_42 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_42 <= _GEN_111;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_43 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_43 <= _GEN_112;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_44 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_44 <= _GEN_113;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_45 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_45 <= _GEN_114;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_46 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_46 <= _GEN_115;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_47 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_47 <= _GEN_116;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_48 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_48 <= _GEN_117;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_49 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_49 <= _GEN_118;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_50 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_50 <= _GEN_119;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_51 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_51 <= _GEN_120;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_52 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_52 <= _GEN_121;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_53 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_53 <= _GEN_122;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_54 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_54 <= _GEN_123;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_55 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_55 <= _GEN_124;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_56 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_56 <= _GEN_125;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_57 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_57 <= _GEN_126;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_58 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_58 <= _GEN_127;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_59 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_59 <= _GEN_128;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_60 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_60 <= _GEN_129;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_61 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_61 <= _GEN_130;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_62 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_62 <= _GEN_131;
        end
      end
    end
    if (io_control == 2'h0) begin // @[WeightedSumModule.scala 40:27]
      buffer_63 <= 18'sh0; // @[WeightedSumModule.scala 42:23]
    end else if (!(io_control == 2'h1)) begin // @[WeightedSumModule.scala 46:33]
      if (!(io_control == 2'h2)) begin // @[WeightedSumModule.scala 63:33]
        if (_T) begin // @[WeightedSumModule.scala 71:33]
          buffer_63 <= _GEN_132;
        end
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      cnt <= 6'h0; // @[Counter.scala 60:40]
    end else if (_T) begin // @[Counter.scala 118:17]
      cnt <= _wrap_value_T_1; // @[Counter.scala 76:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sum = _RAND_0[17:0];
  _RAND_1 = {1{`RANDOM}};
  exp = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  c = _RAND_2[17:0];
  _RAND_3 = {1{`RANDOM}};
  c_exp = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  w1 = _RAND_4[17:0];
  _RAND_5 = {1{`RANDOM}};
  w2 = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  buffer_0 = _RAND_6[17:0];
  _RAND_7 = {1{`RANDOM}};
  buffer_1 = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  buffer_2 = _RAND_8[17:0];
  _RAND_9 = {1{`RANDOM}};
  buffer_3 = _RAND_9[17:0];
  _RAND_10 = {1{`RANDOM}};
  buffer_4 = _RAND_10[17:0];
  _RAND_11 = {1{`RANDOM}};
  buffer_5 = _RAND_11[17:0];
  _RAND_12 = {1{`RANDOM}};
  buffer_6 = _RAND_12[17:0];
  _RAND_13 = {1{`RANDOM}};
  buffer_7 = _RAND_13[17:0];
  _RAND_14 = {1{`RANDOM}};
  buffer_8 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  buffer_9 = _RAND_15[17:0];
  _RAND_16 = {1{`RANDOM}};
  buffer_10 = _RAND_16[17:0];
  _RAND_17 = {1{`RANDOM}};
  buffer_11 = _RAND_17[17:0];
  _RAND_18 = {1{`RANDOM}};
  buffer_12 = _RAND_18[17:0];
  _RAND_19 = {1{`RANDOM}};
  buffer_13 = _RAND_19[17:0];
  _RAND_20 = {1{`RANDOM}};
  buffer_14 = _RAND_20[17:0];
  _RAND_21 = {1{`RANDOM}};
  buffer_15 = _RAND_21[17:0];
  _RAND_22 = {1{`RANDOM}};
  buffer_16 = _RAND_22[17:0];
  _RAND_23 = {1{`RANDOM}};
  buffer_17 = _RAND_23[17:0];
  _RAND_24 = {1{`RANDOM}};
  buffer_18 = _RAND_24[17:0];
  _RAND_25 = {1{`RANDOM}};
  buffer_19 = _RAND_25[17:0];
  _RAND_26 = {1{`RANDOM}};
  buffer_20 = _RAND_26[17:0];
  _RAND_27 = {1{`RANDOM}};
  buffer_21 = _RAND_27[17:0];
  _RAND_28 = {1{`RANDOM}};
  buffer_22 = _RAND_28[17:0];
  _RAND_29 = {1{`RANDOM}};
  buffer_23 = _RAND_29[17:0];
  _RAND_30 = {1{`RANDOM}};
  buffer_24 = _RAND_30[17:0];
  _RAND_31 = {1{`RANDOM}};
  buffer_25 = _RAND_31[17:0];
  _RAND_32 = {1{`RANDOM}};
  buffer_26 = _RAND_32[17:0];
  _RAND_33 = {1{`RANDOM}};
  buffer_27 = _RAND_33[17:0];
  _RAND_34 = {1{`RANDOM}};
  buffer_28 = _RAND_34[17:0];
  _RAND_35 = {1{`RANDOM}};
  buffer_29 = _RAND_35[17:0];
  _RAND_36 = {1{`RANDOM}};
  buffer_30 = _RAND_36[17:0];
  _RAND_37 = {1{`RANDOM}};
  buffer_31 = _RAND_37[17:0];
  _RAND_38 = {1{`RANDOM}};
  buffer_32 = _RAND_38[17:0];
  _RAND_39 = {1{`RANDOM}};
  buffer_33 = _RAND_39[17:0];
  _RAND_40 = {1{`RANDOM}};
  buffer_34 = _RAND_40[17:0];
  _RAND_41 = {1{`RANDOM}};
  buffer_35 = _RAND_41[17:0];
  _RAND_42 = {1{`RANDOM}};
  buffer_36 = _RAND_42[17:0];
  _RAND_43 = {1{`RANDOM}};
  buffer_37 = _RAND_43[17:0];
  _RAND_44 = {1{`RANDOM}};
  buffer_38 = _RAND_44[17:0];
  _RAND_45 = {1{`RANDOM}};
  buffer_39 = _RAND_45[17:0];
  _RAND_46 = {1{`RANDOM}};
  buffer_40 = _RAND_46[17:0];
  _RAND_47 = {1{`RANDOM}};
  buffer_41 = _RAND_47[17:0];
  _RAND_48 = {1{`RANDOM}};
  buffer_42 = _RAND_48[17:0];
  _RAND_49 = {1{`RANDOM}};
  buffer_43 = _RAND_49[17:0];
  _RAND_50 = {1{`RANDOM}};
  buffer_44 = _RAND_50[17:0];
  _RAND_51 = {1{`RANDOM}};
  buffer_45 = _RAND_51[17:0];
  _RAND_52 = {1{`RANDOM}};
  buffer_46 = _RAND_52[17:0];
  _RAND_53 = {1{`RANDOM}};
  buffer_47 = _RAND_53[17:0];
  _RAND_54 = {1{`RANDOM}};
  buffer_48 = _RAND_54[17:0];
  _RAND_55 = {1{`RANDOM}};
  buffer_49 = _RAND_55[17:0];
  _RAND_56 = {1{`RANDOM}};
  buffer_50 = _RAND_56[17:0];
  _RAND_57 = {1{`RANDOM}};
  buffer_51 = _RAND_57[17:0];
  _RAND_58 = {1{`RANDOM}};
  buffer_52 = _RAND_58[17:0];
  _RAND_59 = {1{`RANDOM}};
  buffer_53 = _RAND_59[17:0];
  _RAND_60 = {1{`RANDOM}};
  buffer_54 = _RAND_60[17:0];
  _RAND_61 = {1{`RANDOM}};
  buffer_55 = _RAND_61[17:0];
  _RAND_62 = {1{`RANDOM}};
  buffer_56 = _RAND_62[17:0];
  _RAND_63 = {1{`RANDOM}};
  buffer_57 = _RAND_63[17:0];
  _RAND_64 = {1{`RANDOM}};
  buffer_58 = _RAND_64[17:0];
  _RAND_65 = {1{`RANDOM}};
  buffer_59 = _RAND_65[17:0];
  _RAND_66 = {1{`RANDOM}};
  buffer_60 = _RAND_66[17:0];
  _RAND_67 = {1{`RANDOM}};
  buffer_61 = _RAND_67[17:0];
  _RAND_68 = {1{`RANDOM}};
  buffer_62 = _RAND_68[17:0];
  _RAND_69 = {1{`RANDOM}};
  buffer_63 = _RAND_69[17:0];
  _RAND_70 = {1{`RANDOM}};
  cnt = _RAND_70[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PEArray(
  input         clock,
  input         reset,
  input  [8:0]  io_kv_ports_0,
  input  [8:0]  io_kv_ports_1,
  input  [8:0]  io_kv_ports_2,
  input  [8:0]  io_kv_ports_3,
  input  [8:0]  io_kv_ports_4,
  input  [8:0]  io_kv_ports_5,
  input  [8:0]  io_kv_ports_6,
  input  [8:0]  io_kv_ports_7,
  input  [8:0]  io_kv_ports_8,
  input  [8:0]  io_kv_ports_9,
  input  [8:0]  io_kv_ports_10,
  input  [8:0]  io_kv_ports_11,
  input  [8:0]  io_kv_ports_12,
  input  [8:0]  io_kv_ports_13,
  input  [8:0]  io_kv_ports_14,
  input  [8:0]  io_kv_ports_15,
  input  [8:0]  io_kv_ports_16,
  input  [8:0]  io_kv_ports_17,
  input  [8:0]  io_kv_ports_18,
  input  [8:0]  io_kv_ports_19,
  input  [8:0]  io_kv_ports_20,
  input  [8:0]  io_kv_ports_21,
  input  [8:0]  io_kv_ports_22,
  input  [8:0]  io_kv_ports_23,
  input  [8:0]  io_kv_ports_24,
  input  [8:0]  io_kv_ports_25,
  input  [8:0]  io_kv_ports_26,
  input  [8:0]  io_kv_ports_27,
  input  [8:0]  io_kv_ports_28,
  input  [8:0]  io_kv_ports_29,
  input  [8:0]  io_kv_ports_30,
  input  [8:0]  io_kv_ports_31,
  input  [8:0]  io_kv_ports_32,
  input  [8:0]  io_kv_ports_33,
  input  [8:0]  io_kv_ports_34,
  input  [8:0]  io_kv_ports_35,
  input  [8:0]  io_kv_ports_36,
  input  [8:0]  io_kv_ports_37,
  input  [8:0]  io_kv_ports_38,
  input  [8:0]  io_kv_ports_39,
  input  [8:0]  io_kv_ports_40,
  input  [8:0]  io_kv_ports_41,
  input  [8:0]  io_kv_ports_42,
  input  [8:0]  io_kv_ports_43,
  input  [8:0]  io_kv_ports_44,
  input  [8:0]  io_kv_ports_45,
  input  [8:0]  io_kv_ports_46,
  input  [8:0]  io_kv_ports_47,
  input  [8:0]  io_kv_ports_48,
  input  [8:0]  io_kv_ports_49,
  input  [8:0]  io_kv_ports_50,
  input  [8:0]  io_kv_ports_51,
  input  [8:0]  io_kv_ports_52,
  input  [8:0]  io_kv_ports_53,
  input  [8:0]  io_kv_ports_54,
  input  [8:0]  io_kv_ports_55,
  input  [8:0]  io_kv_ports_56,
  input  [8:0]  io_kv_ports_57,
  input  [8:0]  io_kv_ports_58,
  input  [8:0]  io_kv_ports_59,
  input  [8:0]  io_kv_ports_60,
  input  [8:0]  io_kv_ports_61,
  input  [8:0]  io_kv_ports_62,
  input  [8:0]  io_kv_ports_63,
  input  [8:0]  io_q_ports_0,
  input  [8:0]  io_q_ports_1,
  input  [8:0]  io_q_ports_2,
  input  [8:0]  io_q_ports_3,
  input  [8:0]  io_q_ports_4,
  input  [8:0]  io_q_ports_5,
  input  [8:0]  io_q_ports_6,
  input  [8:0]  io_q_ports_7,
  input  [8:0]  io_q_ports_8,
  input  [8:0]  io_q_ports_9,
  input  [8:0]  io_q_ports_10,
  input  [8:0]  io_q_ports_11,
  input  [8:0]  io_q_ports_12,
  input  [8:0]  io_q_ports_13,
  input  [8:0]  io_q_ports_14,
  input  [8:0]  io_q_ports_15,
  input  [8:0]  io_q_ports_16,
  input  [8:0]  io_q_ports_17,
  input  [8:0]  io_q_ports_18,
  input  [8:0]  io_q_ports_19,
  input  [8:0]  io_q_ports_20,
  input  [8:0]  io_q_ports_21,
  input  [8:0]  io_q_ports_22,
  input  [8:0]  io_q_ports_23,
  input  [8:0]  io_q_ports_24,
  input  [8:0]  io_q_ports_25,
  input  [8:0]  io_q_ports_26,
  input  [8:0]  io_q_ports_27,
  input  [8:0]  io_q_ports_28,
  input  [8:0]  io_q_ports_29,
  input  [8:0]  io_q_ports_30,
  input  [8:0]  io_q_ports_31,
  input  [8:0]  io_q_ports_32,
  input  [2:0]  io_stage_ports_0,
  input  [2:0]  io_stage_ports_1,
  input  [2:0]  io_stage_ports_2,
  input  [2:0]  io_stage_ports_3,
  input  [2:0]  io_stage_ports_4,
  input  [2:0]  io_stage_ports_5,
  input  [2:0]  io_stage_ports_6,
  input  [2:0]  io_stage_ports_7,
  input  [2:0]  io_stage_ports_8,
  input  [2:0]  io_stage_ports_9,
  input  [2:0]  io_stage_ports_10,
  input  [2:0]  io_stage_ports_11,
  input  [2:0]  io_stage_ports_12,
  input  [2:0]  io_stage_ports_13,
  input  [2:0]  io_stage_ports_14,
  input  [2:0]  io_stage_ports_15,
  input  [2:0]  io_stage_ports_16,
  input  [2:0]  io_stage_ports_17,
  input  [2:0]  io_stage_ports_18,
  input  [2:0]  io_stage_ports_19,
  input  [2:0]  io_stage_ports_20,
  input  [2:0]  io_stage_ports_21,
  input  [2:0]  io_stage_ports_22,
  input  [2:0]  io_stage_ports_23,
  input  [2:0]  io_stage_ports_24,
  input  [2:0]  io_stage_ports_25,
  input  [2:0]  io_stage_ports_26,
  input  [2:0]  io_stage_ports_27,
  input  [2:0]  io_stage_ports_28,
  input  [2:0]  io_stage_ports_29,
  input  [2:0]  io_stage_ports_30,
  input  [2:0]  io_stage_ports_31,
  input  [2:0]  io_stage_ports_32,
  input  [1:0]  io_weight_control,
  output [17:0] io_out_ports_0,
  output [17:0] io_out_ports_1,
  output [17:0] io_out_ports_2,
  output [17:0] io_out_ports_3,
  output [17:0] io_out_ports_4,
  output [17:0] io_out_ports_5,
  output [17:0] io_out_ports_6,
  output [17:0] io_out_ports_7,
  output [17:0] io_out_ports_8,
  output [17:0] io_out_ports_9,
  output [17:0] io_out_ports_10,
  output [17:0] io_out_ports_11,
  output [17:0] io_out_ports_12,
  output [17:0] io_out_ports_13,
  output [17:0] io_out_ports_14,
  output [17:0] io_out_ports_15,
  output [17:0] io_out_ports_16,
  output [17:0] io_out_ports_17,
  output [17:0] io_out_ports_18,
  output [17:0] io_out_ports_19,
  output [17:0] io_out_ports_20,
  output [17:0] io_out_ports_21,
  output [17:0] io_out_ports_22,
  output [17:0] io_out_ports_23,
  output [17:0] io_out_ports_24,
  output [17:0] io_out_ports_25,
  output [17:0] io_out_ports_26,
  output [17:0] io_out_ports_27,
  output [17:0] io_out_ports_28,
  output [17:0] io_out_ports_29,
  output [17:0] io_out_ports_30,
  output [17:0] io_out_ports_31,
  output [17:0] io_out_ports_32
);
  wire  local_pes_0_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_0_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_0_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_0_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_0_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_0_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_0_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_1_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_1_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_1_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_1_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_1_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_1_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_2_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_2_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_2_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_2_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_2_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_2_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_3_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_3_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_3_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_3_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_3_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_3_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_4_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_4_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_4_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_4_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_4_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_4_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_5_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_5_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_5_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_5_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_5_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_5_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_6_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_6_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_6_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_6_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_6_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_6_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_7_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_7_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_7_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_7_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_7_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_7_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_8_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_8_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_8_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_8_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_8_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_8_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_9_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_9_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_9_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_9_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_9_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_9_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_10_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_10_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_10_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_10_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_10_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_10_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_11_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_11_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_11_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_11_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_11_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_11_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_12_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_12_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_12_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_12_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_12_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_12_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_13_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_13_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_13_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_13_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_13_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_13_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_14_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_14_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_14_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_14_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_14_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_14_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_15_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_15_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_15_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_15_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_15_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_15_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_16_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_16_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_16_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_16_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_16_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_16_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_17_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_17_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_17_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_17_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_17_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_17_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_18_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_18_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_18_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_18_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_18_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_18_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_19_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_19_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_19_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_19_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_19_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_19_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_20_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_20_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_20_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_20_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_20_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_20_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_21_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_21_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_21_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_21_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_21_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_21_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_22_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_22_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_22_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_22_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_22_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_22_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_23_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_23_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_23_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_23_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_23_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_23_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_24_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_24_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_24_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_24_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_24_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_24_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_25_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_25_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_25_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_25_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_25_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_25_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_26_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_26_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_26_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_26_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_26_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_26_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_27_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_27_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_27_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_27_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_27_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_27_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_28_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_28_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_28_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_28_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_28_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_28_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_29_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_29_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_29_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_29_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_29_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_29_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_30_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_30_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_30_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_30_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_30_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_30_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_0_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_0_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_0_io_in_q; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_0_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_0_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_0_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_0_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_0_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_0_io_out_sum; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_0_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_0_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_1_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_1_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_1_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_1_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_1_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_1_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_1_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_1_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_1_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_1_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_1_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_1_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_1_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_1_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_2_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_2_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_2_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_2_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_2_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_2_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_2_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_2_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_2_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_2_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_2_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_2_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_2_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_2_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_3_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_3_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_3_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_3_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_3_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_3_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_3_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_3_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_3_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_3_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_3_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_3_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_3_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_3_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_4_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_4_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_4_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_4_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_4_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_4_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_4_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_4_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_4_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_4_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_4_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_4_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_4_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_4_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_5_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_5_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_5_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_5_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_5_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_5_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_5_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_5_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_5_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_5_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_5_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_5_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_5_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_5_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_6_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_6_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_6_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_6_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_6_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_6_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_6_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_6_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_6_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_6_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_6_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_6_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_6_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_6_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_7_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_7_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_7_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_7_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_7_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_7_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_7_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_7_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_7_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_7_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_7_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_7_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_7_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_7_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_8_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_8_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_8_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_8_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_8_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_8_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_8_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_8_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_8_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_8_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_8_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_8_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_8_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_8_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_9_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_9_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_9_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_9_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_9_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_9_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_9_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_9_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_9_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_9_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_9_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_9_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_9_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_9_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_10_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_10_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_10_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_10_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_10_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_10_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_10_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_10_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_10_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_10_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_10_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_10_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_10_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_10_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_11_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_11_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_11_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_11_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_11_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_11_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_11_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_11_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_11_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_11_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_11_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_11_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_11_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_11_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_12_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_12_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_12_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_12_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_12_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_12_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_12_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_12_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_12_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_12_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_12_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_12_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_12_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_12_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_13_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_13_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_13_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_13_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_13_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_13_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_13_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_13_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_13_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_13_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_13_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_13_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_13_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_13_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_14_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_14_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_14_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_14_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_14_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_14_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_14_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_14_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_14_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_14_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_14_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_14_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_14_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_14_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_15_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_15_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_15_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_15_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_15_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_15_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_15_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_15_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_15_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_15_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_15_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_15_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_15_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_15_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_16_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_16_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_16_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_16_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_16_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_16_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_16_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_16_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_16_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_16_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_16_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_16_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_16_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_16_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_17_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_17_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_17_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_17_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_17_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_17_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_17_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_17_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_17_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_17_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_17_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_17_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_17_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_17_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_18_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_18_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_18_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_18_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_18_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_18_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_18_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_18_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_18_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_18_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_18_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_18_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_18_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_18_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_19_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_19_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_19_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_19_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_19_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_19_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_19_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_19_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_19_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_19_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_19_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_19_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_19_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_19_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_20_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_20_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_20_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_20_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_20_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_20_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_20_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_20_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_20_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_20_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_20_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_20_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_20_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_20_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_21_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_21_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_21_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_21_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_21_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_21_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_21_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_21_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_21_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_21_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_21_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_21_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_21_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_21_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_22_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_22_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_22_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_22_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_22_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_22_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_22_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_22_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_22_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_22_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_22_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_22_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_22_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_22_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_23_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_23_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_23_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_23_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_23_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_23_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_23_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_23_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_23_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_23_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_23_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_23_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_23_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_23_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_24_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_24_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_24_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_24_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_24_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_24_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_24_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_24_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_24_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_24_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_24_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_24_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_24_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_24_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_25_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_25_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_25_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_25_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_25_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_25_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_25_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_25_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_25_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_25_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_25_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_25_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_25_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_25_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_26_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_26_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_26_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_26_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_26_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_26_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_26_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_26_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_26_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_26_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_26_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_26_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_26_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_26_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_27_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_27_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_27_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_27_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_27_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_27_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_27_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_27_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_27_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_27_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_27_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_27_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_27_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_27_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_28_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_28_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_28_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_28_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_28_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_28_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_28_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_28_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_28_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_28_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_28_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_28_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_28_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_28_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_29_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_29_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_29_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_29_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_29_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_29_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_29_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_29_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_29_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_29_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_29_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_29_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_29_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_29_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_30_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_30_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_30_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_30_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_30_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_30_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_30_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_30_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_30_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_30_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_30_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_30_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_30_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_30_io_out_stage; // @[PEArray.scala 23:49]
  wire  local_pes_31_31_clock; // @[PEArray.scala 23:49]
  wire  local_pes_31_31_reset; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_31_io_in_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_31_io_in_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_31_io_in_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_31_io_in_kv; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_31_io_in_inv_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_31_io_in_inv_sum; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_31_io_in_stage; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_31_io_out_q; // @[PEArray.scala 23:49]
  wire [17:0] local_pes_31_31_io_out_sum; // @[PEArray.scala 23:49]
  wire [4:0] local_pes_31_31_io_out_sum_exp; // @[PEArray.scala 23:49]
  wire [8:0] local_pes_31_31_io_out_kv; // @[PEArray.scala 23:49]
  wire [2:0] local_pes_31_31_io_out_stage; // @[PEArray.scala 23:49]
  wire  global_col_pes_0_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_0_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_0_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_0_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_0_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_0_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_0_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_0_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_0_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_0_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_0_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_0_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_0_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_0_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_1_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_1_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_1_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_1_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_1_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_1_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_1_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_1_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_1_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_1_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_1_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_1_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_1_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_1_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_2_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_2_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_2_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_2_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_2_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_2_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_2_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_2_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_2_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_2_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_2_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_2_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_2_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_2_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_3_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_3_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_3_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_3_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_3_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_3_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_3_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_3_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_3_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_3_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_3_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_3_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_3_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_3_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_4_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_4_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_4_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_4_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_4_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_4_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_4_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_4_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_4_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_4_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_4_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_4_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_4_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_4_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_5_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_5_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_5_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_5_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_5_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_5_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_5_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_5_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_5_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_5_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_5_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_5_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_5_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_5_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_6_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_6_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_6_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_6_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_6_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_6_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_6_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_6_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_6_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_6_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_6_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_6_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_6_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_6_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_7_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_7_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_7_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_7_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_7_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_7_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_7_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_7_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_7_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_7_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_7_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_7_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_7_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_7_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_8_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_8_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_8_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_8_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_8_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_8_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_8_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_8_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_8_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_8_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_8_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_8_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_8_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_8_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_9_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_9_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_9_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_9_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_9_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_9_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_9_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_9_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_9_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_9_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_9_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_9_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_9_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_9_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_10_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_10_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_10_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_10_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_10_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_10_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_10_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_10_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_10_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_10_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_10_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_10_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_10_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_10_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_11_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_11_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_11_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_11_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_11_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_11_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_11_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_11_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_11_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_11_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_11_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_11_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_11_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_11_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_12_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_12_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_12_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_12_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_12_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_12_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_12_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_12_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_12_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_12_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_12_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_12_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_12_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_12_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_13_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_13_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_13_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_13_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_13_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_13_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_13_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_13_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_13_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_13_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_13_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_13_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_13_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_13_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_14_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_14_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_14_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_14_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_14_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_14_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_14_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_14_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_14_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_14_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_14_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_14_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_14_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_14_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_15_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_15_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_15_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_15_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_15_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_15_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_15_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_15_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_15_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_15_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_15_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_15_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_15_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_15_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_16_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_16_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_16_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_16_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_16_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_16_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_16_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_16_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_16_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_16_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_16_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_16_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_16_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_16_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_17_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_17_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_17_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_17_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_17_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_17_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_17_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_17_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_17_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_17_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_17_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_17_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_17_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_17_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_18_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_18_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_18_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_18_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_18_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_18_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_18_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_18_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_18_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_18_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_18_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_18_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_18_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_18_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_19_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_19_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_19_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_19_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_19_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_19_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_19_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_19_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_19_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_19_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_19_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_19_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_19_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_19_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_20_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_20_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_20_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_20_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_20_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_20_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_20_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_20_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_20_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_20_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_20_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_20_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_20_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_20_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_21_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_21_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_21_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_21_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_21_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_21_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_21_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_21_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_21_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_21_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_21_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_21_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_21_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_21_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_22_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_22_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_22_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_22_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_22_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_22_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_22_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_22_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_22_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_22_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_22_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_22_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_22_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_22_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_23_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_23_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_23_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_23_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_23_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_23_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_23_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_23_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_23_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_23_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_23_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_23_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_23_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_23_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_24_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_24_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_24_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_24_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_24_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_24_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_24_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_24_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_24_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_24_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_24_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_24_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_24_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_24_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_25_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_25_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_25_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_25_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_25_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_25_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_25_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_25_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_25_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_25_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_25_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_25_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_25_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_25_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_26_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_26_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_26_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_26_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_26_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_26_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_26_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_26_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_26_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_26_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_26_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_26_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_26_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_26_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_27_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_27_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_27_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_27_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_27_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_27_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_27_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_27_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_27_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_27_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_27_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_27_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_27_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_27_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_28_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_28_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_28_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_28_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_28_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_28_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_28_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_28_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_28_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_28_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_28_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_28_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_28_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_28_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_29_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_29_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_29_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_29_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_29_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_29_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_29_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_29_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_29_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_29_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_29_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_29_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_29_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_29_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_30_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_30_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_30_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_30_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_30_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_30_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_30_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_30_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_30_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_30_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_30_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_30_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_30_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_30_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_col_pes_31_0_clock; // @[PEArray.scala 26:50]
  wire  global_col_pes_31_0_reset; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_31_0_io_in_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_31_0_io_in_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_31_0_io_in_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_31_0_io_in_kv; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_31_0_io_in_inv_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_31_0_io_in_inv_sum; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_31_0_io_in_stage; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_31_0_io_out_q; // @[PEArray.scala 26:50]
  wire [17:0] global_col_pes_31_0_io_out_sum; // @[PEArray.scala 26:50]
  wire [4:0] global_col_pes_31_0_io_out_sum_exp; // @[PEArray.scala 26:50]
  wire [8:0] global_col_pes_31_0_io_out_kv; // @[PEArray.scala 26:50]
  wire [2:0] global_col_pes_31_0_io_out_stage; // @[PEArray.scala 26:50]
  wire  global_row_pes_0_0_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_0_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_0_io_in_q; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_0_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_0_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_0_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_0_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_0_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_0_io_out_sum; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_0_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_0_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_1_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_1_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_1_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_1_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_1_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_1_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_1_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_1_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_1_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_1_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_1_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_1_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_1_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_1_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_2_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_2_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_2_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_2_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_2_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_2_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_2_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_2_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_2_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_2_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_2_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_2_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_2_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_2_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_3_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_3_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_3_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_3_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_3_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_3_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_3_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_3_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_3_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_3_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_3_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_3_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_3_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_3_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_4_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_4_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_4_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_4_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_4_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_4_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_4_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_4_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_4_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_4_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_4_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_4_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_4_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_4_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_5_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_5_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_5_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_5_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_5_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_5_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_5_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_5_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_5_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_5_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_5_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_5_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_5_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_5_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_6_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_6_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_6_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_6_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_6_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_6_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_6_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_6_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_6_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_6_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_6_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_6_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_6_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_6_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_7_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_7_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_7_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_7_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_7_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_7_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_7_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_7_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_7_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_7_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_7_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_7_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_7_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_7_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_8_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_8_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_8_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_8_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_8_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_8_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_8_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_8_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_8_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_8_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_8_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_8_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_8_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_8_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_9_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_9_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_9_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_9_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_9_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_9_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_9_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_9_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_9_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_9_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_9_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_9_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_9_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_9_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_10_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_10_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_10_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_10_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_10_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_10_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_10_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_10_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_10_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_10_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_10_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_10_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_10_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_10_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_11_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_11_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_11_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_11_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_11_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_11_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_11_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_11_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_11_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_11_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_11_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_11_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_11_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_11_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_12_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_12_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_12_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_12_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_12_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_12_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_12_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_12_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_12_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_12_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_12_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_12_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_12_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_12_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_13_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_13_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_13_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_13_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_13_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_13_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_13_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_13_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_13_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_13_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_13_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_13_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_13_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_13_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_14_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_14_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_14_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_14_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_14_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_14_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_14_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_14_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_14_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_14_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_14_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_14_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_14_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_14_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_15_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_15_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_15_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_15_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_15_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_15_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_15_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_15_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_15_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_15_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_15_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_15_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_15_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_15_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_16_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_16_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_16_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_16_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_16_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_16_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_16_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_16_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_16_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_16_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_16_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_16_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_16_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_16_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_17_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_17_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_17_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_17_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_17_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_17_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_17_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_17_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_17_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_17_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_17_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_17_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_17_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_17_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_18_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_18_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_18_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_18_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_18_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_18_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_18_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_18_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_18_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_18_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_18_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_18_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_18_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_18_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_19_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_19_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_19_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_19_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_19_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_19_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_19_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_19_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_19_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_19_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_19_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_19_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_19_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_19_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_20_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_20_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_20_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_20_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_20_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_20_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_20_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_20_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_20_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_20_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_20_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_20_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_20_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_20_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_21_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_21_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_21_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_21_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_21_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_21_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_21_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_21_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_21_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_21_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_21_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_21_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_21_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_21_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_22_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_22_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_22_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_22_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_22_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_22_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_22_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_22_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_22_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_22_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_22_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_22_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_22_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_22_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_23_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_23_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_23_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_23_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_23_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_23_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_23_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_23_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_23_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_23_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_23_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_23_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_23_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_23_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_24_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_24_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_24_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_24_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_24_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_24_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_24_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_24_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_24_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_24_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_24_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_24_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_24_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_24_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_25_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_25_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_25_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_25_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_25_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_25_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_25_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_25_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_25_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_25_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_25_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_25_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_25_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_25_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_26_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_26_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_26_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_26_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_26_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_26_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_26_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_26_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_26_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_26_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_26_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_26_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_26_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_26_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_27_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_27_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_27_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_27_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_27_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_27_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_27_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_27_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_27_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_27_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_27_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_27_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_27_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_27_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_28_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_28_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_28_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_28_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_28_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_28_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_28_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_28_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_28_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_28_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_28_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_28_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_28_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_28_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_29_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_29_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_29_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_29_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_29_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_29_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_29_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_29_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_29_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_29_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_29_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_29_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_29_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_29_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_30_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_30_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_30_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_30_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_30_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_30_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_30_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_30_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_30_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_30_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_30_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_30_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_30_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_30_io_out_stage; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_31_clock; // @[PEArray.scala 29:49]
  wire  global_row_pes_0_31_reset; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_31_io_in_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_31_io_in_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_31_io_in_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_31_io_in_kv; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_31_io_in_inv_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_31_io_in_inv_sum; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_31_io_in_stage; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_31_io_out_q; // @[PEArray.scala 29:49]
  wire [17:0] global_row_pes_0_31_io_out_sum; // @[PEArray.scala 29:49]
  wire [4:0] global_row_pes_0_31_io_out_sum_exp; // @[PEArray.scala 29:49]
  wire [8:0] global_row_pes_0_31_io_out_kv; // @[PEArray.scala 29:49]
  wire [2:0] global_row_pes_0_31_io_out_stage; // @[PEArray.scala 29:49]
  wire [17:0] inv_modules_0_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_0_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_0_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_1_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_1_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_1_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_2_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_2_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_2_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_3_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_3_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_3_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_4_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_4_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_4_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_5_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_5_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_5_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_6_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_6_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_6_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_7_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_7_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_7_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_8_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_8_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_8_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_9_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_9_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_9_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_10_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_10_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_10_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_11_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_11_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_11_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_12_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_12_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_12_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_13_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_13_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_13_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_14_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_14_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_14_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_15_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_15_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_15_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_16_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_16_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_16_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_17_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_17_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_17_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_18_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_18_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_18_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_19_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_19_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_19_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_20_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_20_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_20_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_21_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_21_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_21_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_22_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_22_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_22_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_23_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_23_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_23_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_24_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_24_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_24_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_25_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_25_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_25_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_26_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_26_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_26_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_27_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_27_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_27_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_28_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_28_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_28_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_29_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_29_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_29_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_30_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_30_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_30_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_31_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_31_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_31_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire [17:0] inv_modules_32_io_in_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_32_io_in_exp; // @[PEArray.scala 31:73]
  wire [8:0] inv_modules_32_io_out_inv_sum; // @[PEArray.scala 31:73]
  wire [4:0] inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 31:73]
  wire  weighted_sum_modules_0_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_0_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_0_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_0_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_0_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_0_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_1_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_1_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_1_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_1_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_1_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_1_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_2_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_2_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_2_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_2_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_2_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_2_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_3_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_3_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_3_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_3_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_3_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_3_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_4_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_4_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_4_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_4_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_4_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_4_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_5_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_5_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_5_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_5_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_5_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_5_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_6_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_6_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_6_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_6_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_6_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_6_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_7_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_7_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_7_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_7_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_7_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_7_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_8_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_8_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_8_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_8_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_8_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_8_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_9_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_9_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_9_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_9_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_9_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_9_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_10_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_10_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_10_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_10_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_10_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_10_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_11_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_11_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_11_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_11_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_11_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_11_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_12_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_12_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_12_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_12_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_12_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_12_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_13_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_13_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_13_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_13_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_13_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_13_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_14_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_14_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_14_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_14_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_14_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_14_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_15_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_15_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_15_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_15_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_15_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_15_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_16_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_16_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_16_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_16_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_16_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_16_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_17_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_17_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_17_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_17_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_17_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_17_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_18_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_18_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_18_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_18_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_18_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_18_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_19_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_19_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_19_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_19_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_19_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_19_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_20_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_20_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_20_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_20_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_20_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_20_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_21_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_21_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_21_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_21_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_21_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_21_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_22_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_22_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_22_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_22_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_22_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_22_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_23_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_23_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_23_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_23_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_23_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_23_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_24_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_24_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_24_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_24_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_24_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_24_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_25_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_25_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_25_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_25_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_25_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_25_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_26_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_26_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_26_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_26_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_26_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_26_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_27_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_27_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_27_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_27_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_27_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_27_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_28_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_28_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_28_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_28_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_28_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_28_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_29_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_29_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_29_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_29_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_29_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_29_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_30_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_30_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_30_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_30_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_30_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_30_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_31_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_31_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_31_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_31_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_31_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_31_io_out_port; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_32_clock; // @[PEArray.scala 33:82]
  wire  weighted_sum_modules_32_reset; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_32_io_in_sum; // @[PEArray.scala 33:82]
  wire [4:0] weighted_sum_modules_32_io_in_exp; // @[PEArray.scala 33:82]
  wire [1:0] weighted_sum_modules_32_io_control; // @[PEArray.scala 33:82]
  wire [17:0] weighted_sum_modules_32_io_out_port; // @[PEArray.scala 33:82]
  wire [11:0] _GEN_0 = {$signed(inv_modules_0_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_64 = {$signed(inv_modules_1_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_128 = {$signed(inv_modules_2_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_192 = {$signed(inv_modules_3_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_256 = {$signed(inv_modules_4_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_320 = {$signed(inv_modules_5_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_384 = {$signed(inv_modules_6_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_448 = {$signed(inv_modules_7_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_512 = {$signed(inv_modules_8_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_576 = {$signed(inv_modules_9_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_640 = {$signed(inv_modules_10_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_704 = {$signed(inv_modules_11_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_768 = {$signed(inv_modules_12_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_832 = {$signed(inv_modules_13_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_896 = {$signed(inv_modules_14_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_960 = {$signed(inv_modules_15_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1024 = {$signed(inv_modules_16_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1088 = {$signed(inv_modules_17_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1152 = {$signed(inv_modules_18_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1216 = {$signed(inv_modules_19_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1280 = {$signed(inv_modules_20_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1344 = {$signed(inv_modules_21_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1408 = {$signed(inv_modules_22_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1472 = {$signed(inv_modules_23_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1536 = {$signed(inv_modules_24_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1600 = {$signed(inv_modules_25_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1664 = {$signed(inv_modules_26_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1728 = {$signed(inv_modules_27_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1792 = {$signed(inv_modules_28_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1856 = {$signed(inv_modules_29_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1920 = {$signed(inv_modules_30_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_1984 = {$signed(inv_modules_31_io_out_inv_sum), 3'h0}; // @[PEArray.scala 55:43]
  wire [11:0] _GEN_2112 = {$signed(inv_modules_32_io_out_inv_sum), 3'h0}; // @[PEArray.scala 79:48]
  PE local_pes_0_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_0_clock),
    .reset(local_pes_0_0_reset),
    .io_in_q(local_pes_0_0_io_in_q),
    .io_in_kv(local_pes_0_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_0_io_in_inv_sum),
    .io_in_stage(local_pes_0_0_io_in_stage),
    .io_out_q(local_pes_0_0_io_out_q),
    .io_out_sum(local_pes_0_0_io_out_sum),
    .io_out_kv(local_pes_0_0_io_out_kv),
    .io_out_stage(local_pes_0_0_io_out_stage)
  );
  PE_1 local_pes_0_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_1_clock),
    .reset(local_pes_0_1_reset),
    .io_in_q(local_pes_0_1_io_in_q),
    .io_in_sum(local_pes_0_1_io_in_sum),
    .io_in_sum_exp(local_pes_0_1_io_in_sum_exp),
    .io_in_kv(local_pes_0_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_1_io_in_inv_sum),
    .io_in_stage(local_pes_0_1_io_in_stage),
    .io_out_q(local_pes_0_1_io_out_q),
    .io_out_sum(local_pes_0_1_io_out_sum),
    .io_out_sum_exp(local_pes_0_1_io_out_sum_exp),
    .io_out_kv(local_pes_0_1_io_out_kv),
    .io_out_stage(local_pes_0_1_io_out_stage)
  );
  PE_1 local_pes_0_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_2_clock),
    .reset(local_pes_0_2_reset),
    .io_in_q(local_pes_0_2_io_in_q),
    .io_in_sum(local_pes_0_2_io_in_sum),
    .io_in_sum_exp(local_pes_0_2_io_in_sum_exp),
    .io_in_kv(local_pes_0_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_2_io_in_inv_sum),
    .io_in_stage(local_pes_0_2_io_in_stage),
    .io_out_q(local_pes_0_2_io_out_q),
    .io_out_sum(local_pes_0_2_io_out_sum),
    .io_out_sum_exp(local_pes_0_2_io_out_sum_exp),
    .io_out_kv(local_pes_0_2_io_out_kv),
    .io_out_stage(local_pes_0_2_io_out_stage)
  );
  PE_1 local_pes_0_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_3_clock),
    .reset(local_pes_0_3_reset),
    .io_in_q(local_pes_0_3_io_in_q),
    .io_in_sum(local_pes_0_3_io_in_sum),
    .io_in_sum_exp(local_pes_0_3_io_in_sum_exp),
    .io_in_kv(local_pes_0_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_3_io_in_inv_sum),
    .io_in_stage(local_pes_0_3_io_in_stage),
    .io_out_q(local_pes_0_3_io_out_q),
    .io_out_sum(local_pes_0_3_io_out_sum),
    .io_out_sum_exp(local_pes_0_3_io_out_sum_exp),
    .io_out_kv(local_pes_0_3_io_out_kv),
    .io_out_stage(local_pes_0_3_io_out_stage)
  );
  PE_1 local_pes_0_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_4_clock),
    .reset(local_pes_0_4_reset),
    .io_in_q(local_pes_0_4_io_in_q),
    .io_in_sum(local_pes_0_4_io_in_sum),
    .io_in_sum_exp(local_pes_0_4_io_in_sum_exp),
    .io_in_kv(local_pes_0_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_4_io_in_inv_sum),
    .io_in_stage(local_pes_0_4_io_in_stage),
    .io_out_q(local_pes_0_4_io_out_q),
    .io_out_sum(local_pes_0_4_io_out_sum),
    .io_out_sum_exp(local_pes_0_4_io_out_sum_exp),
    .io_out_kv(local_pes_0_4_io_out_kv),
    .io_out_stage(local_pes_0_4_io_out_stage)
  );
  PE_1 local_pes_0_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_5_clock),
    .reset(local_pes_0_5_reset),
    .io_in_q(local_pes_0_5_io_in_q),
    .io_in_sum(local_pes_0_5_io_in_sum),
    .io_in_sum_exp(local_pes_0_5_io_in_sum_exp),
    .io_in_kv(local_pes_0_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_5_io_in_inv_sum),
    .io_in_stage(local_pes_0_5_io_in_stage),
    .io_out_q(local_pes_0_5_io_out_q),
    .io_out_sum(local_pes_0_5_io_out_sum),
    .io_out_sum_exp(local_pes_0_5_io_out_sum_exp),
    .io_out_kv(local_pes_0_5_io_out_kv),
    .io_out_stage(local_pes_0_5_io_out_stage)
  );
  PE_1 local_pes_0_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_6_clock),
    .reset(local_pes_0_6_reset),
    .io_in_q(local_pes_0_6_io_in_q),
    .io_in_sum(local_pes_0_6_io_in_sum),
    .io_in_sum_exp(local_pes_0_6_io_in_sum_exp),
    .io_in_kv(local_pes_0_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_6_io_in_inv_sum),
    .io_in_stage(local_pes_0_6_io_in_stage),
    .io_out_q(local_pes_0_6_io_out_q),
    .io_out_sum(local_pes_0_6_io_out_sum),
    .io_out_sum_exp(local_pes_0_6_io_out_sum_exp),
    .io_out_kv(local_pes_0_6_io_out_kv),
    .io_out_stage(local_pes_0_6_io_out_stage)
  );
  PE_1 local_pes_0_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_7_clock),
    .reset(local_pes_0_7_reset),
    .io_in_q(local_pes_0_7_io_in_q),
    .io_in_sum(local_pes_0_7_io_in_sum),
    .io_in_sum_exp(local_pes_0_7_io_in_sum_exp),
    .io_in_kv(local_pes_0_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_7_io_in_inv_sum),
    .io_in_stage(local_pes_0_7_io_in_stage),
    .io_out_q(local_pes_0_7_io_out_q),
    .io_out_sum(local_pes_0_7_io_out_sum),
    .io_out_sum_exp(local_pes_0_7_io_out_sum_exp),
    .io_out_kv(local_pes_0_7_io_out_kv),
    .io_out_stage(local_pes_0_7_io_out_stage)
  );
  PE_1 local_pes_0_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_8_clock),
    .reset(local_pes_0_8_reset),
    .io_in_q(local_pes_0_8_io_in_q),
    .io_in_sum(local_pes_0_8_io_in_sum),
    .io_in_sum_exp(local_pes_0_8_io_in_sum_exp),
    .io_in_kv(local_pes_0_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_8_io_in_inv_sum),
    .io_in_stage(local_pes_0_8_io_in_stage),
    .io_out_q(local_pes_0_8_io_out_q),
    .io_out_sum(local_pes_0_8_io_out_sum),
    .io_out_sum_exp(local_pes_0_8_io_out_sum_exp),
    .io_out_kv(local_pes_0_8_io_out_kv),
    .io_out_stage(local_pes_0_8_io_out_stage)
  );
  PE_1 local_pes_0_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_9_clock),
    .reset(local_pes_0_9_reset),
    .io_in_q(local_pes_0_9_io_in_q),
    .io_in_sum(local_pes_0_9_io_in_sum),
    .io_in_sum_exp(local_pes_0_9_io_in_sum_exp),
    .io_in_kv(local_pes_0_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_9_io_in_inv_sum),
    .io_in_stage(local_pes_0_9_io_in_stage),
    .io_out_q(local_pes_0_9_io_out_q),
    .io_out_sum(local_pes_0_9_io_out_sum),
    .io_out_sum_exp(local_pes_0_9_io_out_sum_exp),
    .io_out_kv(local_pes_0_9_io_out_kv),
    .io_out_stage(local_pes_0_9_io_out_stage)
  );
  PE_1 local_pes_0_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_10_clock),
    .reset(local_pes_0_10_reset),
    .io_in_q(local_pes_0_10_io_in_q),
    .io_in_sum(local_pes_0_10_io_in_sum),
    .io_in_sum_exp(local_pes_0_10_io_in_sum_exp),
    .io_in_kv(local_pes_0_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_10_io_in_inv_sum),
    .io_in_stage(local_pes_0_10_io_in_stage),
    .io_out_q(local_pes_0_10_io_out_q),
    .io_out_sum(local_pes_0_10_io_out_sum),
    .io_out_sum_exp(local_pes_0_10_io_out_sum_exp),
    .io_out_kv(local_pes_0_10_io_out_kv),
    .io_out_stage(local_pes_0_10_io_out_stage)
  );
  PE_1 local_pes_0_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_11_clock),
    .reset(local_pes_0_11_reset),
    .io_in_q(local_pes_0_11_io_in_q),
    .io_in_sum(local_pes_0_11_io_in_sum),
    .io_in_sum_exp(local_pes_0_11_io_in_sum_exp),
    .io_in_kv(local_pes_0_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_11_io_in_inv_sum),
    .io_in_stage(local_pes_0_11_io_in_stage),
    .io_out_q(local_pes_0_11_io_out_q),
    .io_out_sum(local_pes_0_11_io_out_sum),
    .io_out_sum_exp(local_pes_0_11_io_out_sum_exp),
    .io_out_kv(local_pes_0_11_io_out_kv),
    .io_out_stage(local_pes_0_11_io_out_stage)
  );
  PE_1 local_pes_0_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_12_clock),
    .reset(local_pes_0_12_reset),
    .io_in_q(local_pes_0_12_io_in_q),
    .io_in_sum(local_pes_0_12_io_in_sum),
    .io_in_sum_exp(local_pes_0_12_io_in_sum_exp),
    .io_in_kv(local_pes_0_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_12_io_in_inv_sum),
    .io_in_stage(local_pes_0_12_io_in_stage),
    .io_out_q(local_pes_0_12_io_out_q),
    .io_out_sum(local_pes_0_12_io_out_sum),
    .io_out_sum_exp(local_pes_0_12_io_out_sum_exp),
    .io_out_kv(local_pes_0_12_io_out_kv),
    .io_out_stage(local_pes_0_12_io_out_stage)
  );
  PE_1 local_pes_0_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_13_clock),
    .reset(local_pes_0_13_reset),
    .io_in_q(local_pes_0_13_io_in_q),
    .io_in_sum(local_pes_0_13_io_in_sum),
    .io_in_sum_exp(local_pes_0_13_io_in_sum_exp),
    .io_in_kv(local_pes_0_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_13_io_in_inv_sum),
    .io_in_stage(local_pes_0_13_io_in_stage),
    .io_out_q(local_pes_0_13_io_out_q),
    .io_out_sum(local_pes_0_13_io_out_sum),
    .io_out_sum_exp(local_pes_0_13_io_out_sum_exp),
    .io_out_kv(local_pes_0_13_io_out_kv),
    .io_out_stage(local_pes_0_13_io_out_stage)
  );
  PE_1 local_pes_0_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_14_clock),
    .reset(local_pes_0_14_reset),
    .io_in_q(local_pes_0_14_io_in_q),
    .io_in_sum(local_pes_0_14_io_in_sum),
    .io_in_sum_exp(local_pes_0_14_io_in_sum_exp),
    .io_in_kv(local_pes_0_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_14_io_in_inv_sum),
    .io_in_stage(local_pes_0_14_io_in_stage),
    .io_out_q(local_pes_0_14_io_out_q),
    .io_out_sum(local_pes_0_14_io_out_sum),
    .io_out_sum_exp(local_pes_0_14_io_out_sum_exp),
    .io_out_kv(local_pes_0_14_io_out_kv),
    .io_out_stage(local_pes_0_14_io_out_stage)
  );
  PE_1 local_pes_0_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_15_clock),
    .reset(local_pes_0_15_reset),
    .io_in_q(local_pes_0_15_io_in_q),
    .io_in_sum(local_pes_0_15_io_in_sum),
    .io_in_sum_exp(local_pes_0_15_io_in_sum_exp),
    .io_in_kv(local_pes_0_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_15_io_in_inv_sum),
    .io_in_stage(local_pes_0_15_io_in_stage),
    .io_out_q(local_pes_0_15_io_out_q),
    .io_out_sum(local_pes_0_15_io_out_sum),
    .io_out_sum_exp(local_pes_0_15_io_out_sum_exp),
    .io_out_kv(local_pes_0_15_io_out_kv),
    .io_out_stage(local_pes_0_15_io_out_stage)
  );
  PE_1 local_pes_0_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_16_clock),
    .reset(local_pes_0_16_reset),
    .io_in_q(local_pes_0_16_io_in_q),
    .io_in_sum(local_pes_0_16_io_in_sum),
    .io_in_sum_exp(local_pes_0_16_io_in_sum_exp),
    .io_in_kv(local_pes_0_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_16_io_in_inv_sum),
    .io_in_stage(local_pes_0_16_io_in_stage),
    .io_out_q(local_pes_0_16_io_out_q),
    .io_out_sum(local_pes_0_16_io_out_sum),
    .io_out_sum_exp(local_pes_0_16_io_out_sum_exp),
    .io_out_kv(local_pes_0_16_io_out_kv),
    .io_out_stage(local_pes_0_16_io_out_stage)
  );
  PE_1 local_pes_0_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_17_clock),
    .reset(local_pes_0_17_reset),
    .io_in_q(local_pes_0_17_io_in_q),
    .io_in_sum(local_pes_0_17_io_in_sum),
    .io_in_sum_exp(local_pes_0_17_io_in_sum_exp),
    .io_in_kv(local_pes_0_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_17_io_in_inv_sum),
    .io_in_stage(local_pes_0_17_io_in_stage),
    .io_out_q(local_pes_0_17_io_out_q),
    .io_out_sum(local_pes_0_17_io_out_sum),
    .io_out_sum_exp(local_pes_0_17_io_out_sum_exp),
    .io_out_kv(local_pes_0_17_io_out_kv),
    .io_out_stage(local_pes_0_17_io_out_stage)
  );
  PE_1 local_pes_0_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_18_clock),
    .reset(local_pes_0_18_reset),
    .io_in_q(local_pes_0_18_io_in_q),
    .io_in_sum(local_pes_0_18_io_in_sum),
    .io_in_sum_exp(local_pes_0_18_io_in_sum_exp),
    .io_in_kv(local_pes_0_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_18_io_in_inv_sum),
    .io_in_stage(local_pes_0_18_io_in_stage),
    .io_out_q(local_pes_0_18_io_out_q),
    .io_out_sum(local_pes_0_18_io_out_sum),
    .io_out_sum_exp(local_pes_0_18_io_out_sum_exp),
    .io_out_kv(local_pes_0_18_io_out_kv),
    .io_out_stage(local_pes_0_18_io_out_stage)
  );
  PE_1 local_pes_0_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_19_clock),
    .reset(local_pes_0_19_reset),
    .io_in_q(local_pes_0_19_io_in_q),
    .io_in_sum(local_pes_0_19_io_in_sum),
    .io_in_sum_exp(local_pes_0_19_io_in_sum_exp),
    .io_in_kv(local_pes_0_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_19_io_in_inv_sum),
    .io_in_stage(local_pes_0_19_io_in_stage),
    .io_out_q(local_pes_0_19_io_out_q),
    .io_out_sum(local_pes_0_19_io_out_sum),
    .io_out_sum_exp(local_pes_0_19_io_out_sum_exp),
    .io_out_kv(local_pes_0_19_io_out_kv),
    .io_out_stage(local_pes_0_19_io_out_stage)
  );
  PE_1 local_pes_0_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_20_clock),
    .reset(local_pes_0_20_reset),
    .io_in_q(local_pes_0_20_io_in_q),
    .io_in_sum(local_pes_0_20_io_in_sum),
    .io_in_sum_exp(local_pes_0_20_io_in_sum_exp),
    .io_in_kv(local_pes_0_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_20_io_in_inv_sum),
    .io_in_stage(local_pes_0_20_io_in_stage),
    .io_out_q(local_pes_0_20_io_out_q),
    .io_out_sum(local_pes_0_20_io_out_sum),
    .io_out_sum_exp(local_pes_0_20_io_out_sum_exp),
    .io_out_kv(local_pes_0_20_io_out_kv),
    .io_out_stage(local_pes_0_20_io_out_stage)
  );
  PE_1 local_pes_0_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_21_clock),
    .reset(local_pes_0_21_reset),
    .io_in_q(local_pes_0_21_io_in_q),
    .io_in_sum(local_pes_0_21_io_in_sum),
    .io_in_sum_exp(local_pes_0_21_io_in_sum_exp),
    .io_in_kv(local_pes_0_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_21_io_in_inv_sum),
    .io_in_stage(local_pes_0_21_io_in_stage),
    .io_out_q(local_pes_0_21_io_out_q),
    .io_out_sum(local_pes_0_21_io_out_sum),
    .io_out_sum_exp(local_pes_0_21_io_out_sum_exp),
    .io_out_kv(local_pes_0_21_io_out_kv),
    .io_out_stage(local_pes_0_21_io_out_stage)
  );
  PE_1 local_pes_0_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_22_clock),
    .reset(local_pes_0_22_reset),
    .io_in_q(local_pes_0_22_io_in_q),
    .io_in_sum(local_pes_0_22_io_in_sum),
    .io_in_sum_exp(local_pes_0_22_io_in_sum_exp),
    .io_in_kv(local_pes_0_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_22_io_in_inv_sum),
    .io_in_stage(local_pes_0_22_io_in_stage),
    .io_out_q(local_pes_0_22_io_out_q),
    .io_out_sum(local_pes_0_22_io_out_sum),
    .io_out_sum_exp(local_pes_0_22_io_out_sum_exp),
    .io_out_kv(local_pes_0_22_io_out_kv),
    .io_out_stage(local_pes_0_22_io_out_stage)
  );
  PE_1 local_pes_0_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_23_clock),
    .reset(local_pes_0_23_reset),
    .io_in_q(local_pes_0_23_io_in_q),
    .io_in_sum(local_pes_0_23_io_in_sum),
    .io_in_sum_exp(local_pes_0_23_io_in_sum_exp),
    .io_in_kv(local_pes_0_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_23_io_in_inv_sum),
    .io_in_stage(local_pes_0_23_io_in_stage),
    .io_out_q(local_pes_0_23_io_out_q),
    .io_out_sum(local_pes_0_23_io_out_sum),
    .io_out_sum_exp(local_pes_0_23_io_out_sum_exp),
    .io_out_kv(local_pes_0_23_io_out_kv),
    .io_out_stage(local_pes_0_23_io_out_stage)
  );
  PE_1 local_pes_0_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_24_clock),
    .reset(local_pes_0_24_reset),
    .io_in_q(local_pes_0_24_io_in_q),
    .io_in_sum(local_pes_0_24_io_in_sum),
    .io_in_sum_exp(local_pes_0_24_io_in_sum_exp),
    .io_in_kv(local_pes_0_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_24_io_in_inv_sum),
    .io_in_stage(local_pes_0_24_io_in_stage),
    .io_out_q(local_pes_0_24_io_out_q),
    .io_out_sum(local_pes_0_24_io_out_sum),
    .io_out_sum_exp(local_pes_0_24_io_out_sum_exp),
    .io_out_kv(local_pes_0_24_io_out_kv),
    .io_out_stage(local_pes_0_24_io_out_stage)
  );
  PE_1 local_pes_0_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_25_clock),
    .reset(local_pes_0_25_reset),
    .io_in_q(local_pes_0_25_io_in_q),
    .io_in_sum(local_pes_0_25_io_in_sum),
    .io_in_sum_exp(local_pes_0_25_io_in_sum_exp),
    .io_in_kv(local_pes_0_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_25_io_in_inv_sum),
    .io_in_stage(local_pes_0_25_io_in_stage),
    .io_out_q(local_pes_0_25_io_out_q),
    .io_out_sum(local_pes_0_25_io_out_sum),
    .io_out_sum_exp(local_pes_0_25_io_out_sum_exp),
    .io_out_kv(local_pes_0_25_io_out_kv),
    .io_out_stage(local_pes_0_25_io_out_stage)
  );
  PE_1 local_pes_0_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_26_clock),
    .reset(local_pes_0_26_reset),
    .io_in_q(local_pes_0_26_io_in_q),
    .io_in_sum(local_pes_0_26_io_in_sum),
    .io_in_sum_exp(local_pes_0_26_io_in_sum_exp),
    .io_in_kv(local_pes_0_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_26_io_in_inv_sum),
    .io_in_stage(local_pes_0_26_io_in_stage),
    .io_out_q(local_pes_0_26_io_out_q),
    .io_out_sum(local_pes_0_26_io_out_sum),
    .io_out_sum_exp(local_pes_0_26_io_out_sum_exp),
    .io_out_kv(local_pes_0_26_io_out_kv),
    .io_out_stage(local_pes_0_26_io_out_stage)
  );
  PE_1 local_pes_0_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_27_clock),
    .reset(local_pes_0_27_reset),
    .io_in_q(local_pes_0_27_io_in_q),
    .io_in_sum(local_pes_0_27_io_in_sum),
    .io_in_sum_exp(local_pes_0_27_io_in_sum_exp),
    .io_in_kv(local_pes_0_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_27_io_in_inv_sum),
    .io_in_stage(local_pes_0_27_io_in_stage),
    .io_out_q(local_pes_0_27_io_out_q),
    .io_out_sum(local_pes_0_27_io_out_sum),
    .io_out_sum_exp(local_pes_0_27_io_out_sum_exp),
    .io_out_kv(local_pes_0_27_io_out_kv),
    .io_out_stage(local_pes_0_27_io_out_stage)
  );
  PE_1 local_pes_0_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_28_clock),
    .reset(local_pes_0_28_reset),
    .io_in_q(local_pes_0_28_io_in_q),
    .io_in_sum(local_pes_0_28_io_in_sum),
    .io_in_sum_exp(local_pes_0_28_io_in_sum_exp),
    .io_in_kv(local_pes_0_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_28_io_in_inv_sum),
    .io_in_stage(local_pes_0_28_io_in_stage),
    .io_out_q(local_pes_0_28_io_out_q),
    .io_out_sum(local_pes_0_28_io_out_sum),
    .io_out_sum_exp(local_pes_0_28_io_out_sum_exp),
    .io_out_kv(local_pes_0_28_io_out_kv),
    .io_out_stage(local_pes_0_28_io_out_stage)
  );
  PE_1 local_pes_0_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_29_clock),
    .reset(local_pes_0_29_reset),
    .io_in_q(local_pes_0_29_io_in_q),
    .io_in_sum(local_pes_0_29_io_in_sum),
    .io_in_sum_exp(local_pes_0_29_io_in_sum_exp),
    .io_in_kv(local_pes_0_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_29_io_in_inv_sum),
    .io_in_stage(local_pes_0_29_io_in_stage),
    .io_out_q(local_pes_0_29_io_out_q),
    .io_out_sum(local_pes_0_29_io_out_sum),
    .io_out_sum_exp(local_pes_0_29_io_out_sum_exp),
    .io_out_kv(local_pes_0_29_io_out_kv),
    .io_out_stage(local_pes_0_29_io_out_stage)
  );
  PE_1 local_pes_0_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_30_clock),
    .reset(local_pes_0_30_reset),
    .io_in_q(local_pes_0_30_io_in_q),
    .io_in_sum(local_pes_0_30_io_in_sum),
    .io_in_sum_exp(local_pes_0_30_io_in_sum_exp),
    .io_in_kv(local_pes_0_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_30_io_in_inv_sum),
    .io_in_stage(local_pes_0_30_io_in_stage),
    .io_out_q(local_pes_0_30_io_out_q),
    .io_out_sum(local_pes_0_30_io_out_sum),
    .io_out_sum_exp(local_pes_0_30_io_out_sum_exp),
    .io_out_kv(local_pes_0_30_io_out_kv),
    .io_out_stage(local_pes_0_30_io_out_stage)
  );
  PE_1 local_pes_0_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_0_31_clock),
    .reset(local_pes_0_31_reset),
    .io_in_q(local_pes_0_31_io_in_q),
    .io_in_sum(local_pes_0_31_io_in_sum),
    .io_in_sum_exp(local_pes_0_31_io_in_sum_exp),
    .io_in_kv(local_pes_0_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_0_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_0_31_io_in_inv_sum),
    .io_in_stage(local_pes_0_31_io_in_stage),
    .io_out_q(local_pes_0_31_io_out_q),
    .io_out_sum(local_pes_0_31_io_out_sum),
    .io_out_sum_exp(local_pes_0_31_io_out_sum_exp),
    .io_out_kv(local_pes_0_31_io_out_kv),
    .io_out_stage(local_pes_0_31_io_out_stage)
  );
  PE local_pes_1_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_0_clock),
    .reset(local_pes_1_0_reset),
    .io_in_q(local_pes_1_0_io_in_q),
    .io_in_kv(local_pes_1_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_0_io_in_inv_sum),
    .io_in_stage(local_pes_1_0_io_in_stage),
    .io_out_q(local_pes_1_0_io_out_q),
    .io_out_sum(local_pes_1_0_io_out_sum),
    .io_out_kv(local_pes_1_0_io_out_kv),
    .io_out_stage(local_pes_1_0_io_out_stage)
  );
  PE_1 local_pes_1_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_1_clock),
    .reset(local_pes_1_1_reset),
    .io_in_q(local_pes_1_1_io_in_q),
    .io_in_sum(local_pes_1_1_io_in_sum),
    .io_in_sum_exp(local_pes_1_1_io_in_sum_exp),
    .io_in_kv(local_pes_1_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_1_io_in_inv_sum),
    .io_in_stage(local_pes_1_1_io_in_stage),
    .io_out_q(local_pes_1_1_io_out_q),
    .io_out_sum(local_pes_1_1_io_out_sum),
    .io_out_sum_exp(local_pes_1_1_io_out_sum_exp),
    .io_out_kv(local_pes_1_1_io_out_kv),
    .io_out_stage(local_pes_1_1_io_out_stage)
  );
  PE_1 local_pes_1_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_2_clock),
    .reset(local_pes_1_2_reset),
    .io_in_q(local_pes_1_2_io_in_q),
    .io_in_sum(local_pes_1_2_io_in_sum),
    .io_in_sum_exp(local_pes_1_2_io_in_sum_exp),
    .io_in_kv(local_pes_1_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_2_io_in_inv_sum),
    .io_in_stage(local_pes_1_2_io_in_stage),
    .io_out_q(local_pes_1_2_io_out_q),
    .io_out_sum(local_pes_1_2_io_out_sum),
    .io_out_sum_exp(local_pes_1_2_io_out_sum_exp),
    .io_out_kv(local_pes_1_2_io_out_kv),
    .io_out_stage(local_pes_1_2_io_out_stage)
  );
  PE_1 local_pes_1_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_3_clock),
    .reset(local_pes_1_3_reset),
    .io_in_q(local_pes_1_3_io_in_q),
    .io_in_sum(local_pes_1_3_io_in_sum),
    .io_in_sum_exp(local_pes_1_3_io_in_sum_exp),
    .io_in_kv(local_pes_1_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_3_io_in_inv_sum),
    .io_in_stage(local_pes_1_3_io_in_stage),
    .io_out_q(local_pes_1_3_io_out_q),
    .io_out_sum(local_pes_1_3_io_out_sum),
    .io_out_sum_exp(local_pes_1_3_io_out_sum_exp),
    .io_out_kv(local_pes_1_3_io_out_kv),
    .io_out_stage(local_pes_1_3_io_out_stage)
  );
  PE_1 local_pes_1_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_4_clock),
    .reset(local_pes_1_4_reset),
    .io_in_q(local_pes_1_4_io_in_q),
    .io_in_sum(local_pes_1_4_io_in_sum),
    .io_in_sum_exp(local_pes_1_4_io_in_sum_exp),
    .io_in_kv(local_pes_1_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_4_io_in_inv_sum),
    .io_in_stage(local_pes_1_4_io_in_stage),
    .io_out_q(local_pes_1_4_io_out_q),
    .io_out_sum(local_pes_1_4_io_out_sum),
    .io_out_sum_exp(local_pes_1_4_io_out_sum_exp),
    .io_out_kv(local_pes_1_4_io_out_kv),
    .io_out_stage(local_pes_1_4_io_out_stage)
  );
  PE_1 local_pes_1_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_5_clock),
    .reset(local_pes_1_5_reset),
    .io_in_q(local_pes_1_5_io_in_q),
    .io_in_sum(local_pes_1_5_io_in_sum),
    .io_in_sum_exp(local_pes_1_5_io_in_sum_exp),
    .io_in_kv(local_pes_1_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_5_io_in_inv_sum),
    .io_in_stage(local_pes_1_5_io_in_stage),
    .io_out_q(local_pes_1_5_io_out_q),
    .io_out_sum(local_pes_1_5_io_out_sum),
    .io_out_sum_exp(local_pes_1_5_io_out_sum_exp),
    .io_out_kv(local_pes_1_5_io_out_kv),
    .io_out_stage(local_pes_1_5_io_out_stage)
  );
  PE_1 local_pes_1_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_6_clock),
    .reset(local_pes_1_6_reset),
    .io_in_q(local_pes_1_6_io_in_q),
    .io_in_sum(local_pes_1_6_io_in_sum),
    .io_in_sum_exp(local_pes_1_6_io_in_sum_exp),
    .io_in_kv(local_pes_1_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_6_io_in_inv_sum),
    .io_in_stage(local_pes_1_6_io_in_stage),
    .io_out_q(local_pes_1_6_io_out_q),
    .io_out_sum(local_pes_1_6_io_out_sum),
    .io_out_sum_exp(local_pes_1_6_io_out_sum_exp),
    .io_out_kv(local_pes_1_6_io_out_kv),
    .io_out_stage(local_pes_1_6_io_out_stage)
  );
  PE_1 local_pes_1_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_7_clock),
    .reset(local_pes_1_7_reset),
    .io_in_q(local_pes_1_7_io_in_q),
    .io_in_sum(local_pes_1_7_io_in_sum),
    .io_in_sum_exp(local_pes_1_7_io_in_sum_exp),
    .io_in_kv(local_pes_1_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_7_io_in_inv_sum),
    .io_in_stage(local_pes_1_7_io_in_stage),
    .io_out_q(local_pes_1_7_io_out_q),
    .io_out_sum(local_pes_1_7_io_out_sum),
    .io_out_sum_exp(local_pes_1_7_io_out_sum_exp),
    .io_out_kv(local_pes_1_7_io_out_kv),
    .io_out_stage(local_pes_1_7_io_out_stage)
  );
  PE_1 local_pes_1_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_8_clock),
    .reset(local_pes_1_8_reset),
    .io_in_q(local_pes_1_8_io_in_q),
    .io_in_sum(local_pes_1_8_io_in_sum),
    .io_in_sum_exp(local_pes_1_8_io_in_sum_exp),
    .io_in_kv(local_pes_1_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_8_io_in_inv_sum),
    .io_in_stage(local_pes_1_8_io_in_stage),
    .io_out_q(local_pes_1_8_io_out_q),
    .io_out_sum(local_pes_1_8_io_out_sum),
    .io_out_sum_exp(local_pes_1_8_io_out_sum_exp),
    .io_out_kv(local_pes_1_8_io_out_kv),
    .io_out_stage(local_pes_1_8_io_out_stage)
  );
  PE_1 local_pes_1_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_9_clock),
    .reset(local_pes_1_9_reset),
    .io_in_q(local_pes_1_9_io_in_q),
    .io_in_sum(local_pes_1_9_io_in_sum),
    .io_in_sum_exp(local_pes_1_9_io_in_sum_exp),
    .io_in_kv(local_pes_1_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_9_io_in_inv_sum),
    .io_in_stage(local_pes_1_9_io_in_stage),
    .io_out_q(local_pes_1_9_io_out_q),
    .io_out_sum(local_pes_1_9_io_out_sum),
    .io_out_sum_exp(local_pes_1_9_io_out_sum_exp),
    .io_out_kv(local_pes_1_9_io_out_kv),
    .io_out_stage(local_pes_1_9_io_out_stage)
  );
  PE_1 local_pes_1_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_10_clock),
    .reset(local_pes_1_10_reset),
    .io_in_q(local_pes_1_10_io_in_q),
    .io_in_sum(local_pes_1_10_io_in_sum),
    .io_in_sum_exp(local_pes_1_10_io_in_sum_exp),
    .io_in_kv(local_pes_1_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_10_io_in_inv_sum),
    .io_in_stage(local_pes_1_10_io_in_stage),
    .io_out_q(local_pes_1_10_io_out_q),
    .io_out_sum(local_pes_1_10_io_out_sum),
    .io_out_sum_exp(local_pes_1_10_io_out_sum_exp),
    .io_out_kv(local_pes_1_10_io_out_kv),
    .io_out_stage(local_pes_1_10_io_out_stage)
  );
  PE_1 local_pes_1_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_11_clock),
    .reset(local_pes_1_11_reset),
    .io_in_q(local_pes_1_11_io_in_q),
    .io_in_sum(local_pes_1_11_io_in_sum),
    .io_in_sum_exp(local_pes_1_11_io_in_sum_exp),
    .io_in_kv(local_pes_1_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_11_io_in_inv_sum),
    .io_in_stage(local_pes_1_11_io_in_stage),
    .io_out_q(local_pes_1_11_io_out_q),
    .io_out_sum(local_pes_1_11_io_out_sum),
    .io_out_sum_exp(local_pes_1_11_io_out_sum_exp),
    .io_out_kv(local_pes_1_11_io_out_kv),
    .io_out_stage(local_pes_1_11_io_out_stage)
  );
  PE_1 local_pes_1_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_12_clock),
    .reset(local_pes_1_12_reset),
    .io_in_q(local_pes_1_12_io_in_q),
    .io_in_sum(local_pes_1_12_io_in_sum),
    .io_in_sum_exp(local_pes_1_12_io_in_sum_exp),
    .io_in_kv(local_pes_1_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_12_io_in_inv_sum),
    .io_in_stage(local_pes_1_12_io_in_stage),
    .io_out_q(local_pes_1_12_io_out_q),
    .io_out_sum(local_pes_1_12_io_out_sum),
    .io_out_sum_exp(local_pes_1_12_io_out_sum_exp),
    .io_out_kv(local_pes_1_12_io_out_kv),
    .io_out_stage(local_pes_1_12_io_out_stage)
  );
  PE_1 local_pes_1_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_13_clock),
    .reset(local_pes_1_13_reset),
    .io_in_q(local_pes_1_13_io_in_q),
    .io_in_sum(local_pes_1_13_io_in_sum),
    .io_in_sum_exp(local_pes_1_13_io_in_sum_exp),
    .io_in_kv(local_pes_1_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_13_io_in_inv_sum),
    .io_in_stage(local_pes_1_13_io_in_stage),
    .io_out_q(local_pes_1_13_io_out_q),
    .io_out_sum(local_pes_1_13_io_out_sum),
    .io_out_sum_exp(local_pes_1_13_io_out_sum_exp),
    .io_out_kv(local_pes_1_13_io_out_kv),
    .io_out_stage(local_pes_1_13_io_out_stage)
  );
  PE_1 local_pes_1_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_14_clock),
    .reset(local_pes_1_14_reset),
    .io_in_q(local_pes_1_14_io_in_q),
    .io_in_sum(local_pes_1_14_io_in_sum),
    .io_in_sum_exp(local_pes_1_14_io_in_sum_exp),
    .io_in_kv(local_pes_1_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_14_io_in_inv_sum),
    .io_in_stage(local_pes_1_14_io_in_stage),
    .io_out_q(local_pes_1_14_io_out_q),
    .io_out_sum(local_pes_1_14_io_out_sum),
    .io_out_sum_exp(local_pes_1_14_io_out_sum_exp),
    .io_out_kv(local_pes_1_14_io_out_kv),
    .io_out_stage(local_pes_1_14_io_out_stage)
  );
  PE_1 local_pes_1_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_15_clock),
    .reset(local_pes_1_15_reset),
    .io_in_q(local_pes_1_15_io_in_q),
    .io_in_sum(local_pes_1_15_io_in_sum),
    .io_in_sum_exp(local_pes_1_15_io_in_sum_exp),
    .io_in_kv(local_pes_1_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_15_io_in_inv_sum),
    .io_in_stage(local_pes_1_15_io_in_stage),
    .io_out_q(local_pes_1_15_io_out_q),
    .io_out_sum(local_pes_1_15_io_out_sum),
    .io_out_sum_exp(local_pes_1_15_io_out_sum_exp),
    .io_out_kv(local_pes_1_15_io_out_kv),
    .io_out_stage(local_pes_1_15_io_out_stage)
  );
  PE_1 local_pes_1_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_16_clock),
    .reset(local_pes_1_16_reset),
    .io_in_q(local_pes_1_16_io_in_q),
    .io_in_sum(local_pes_1_16_io_in_sum),
    .io_in_sum_exp(local_pes_1_16_io_in_sum_exp),
    .io_in_kv(local_pes_1_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_16_io_in_inv_sum),
    .io_in_stage(local_pes_1_16_io_in_stage),
    .io_out_q(local_pes_1_16_io_out_q),
    .io_out_sum(local_pes_1_16_io_out_sum),
    .io_out_sum_exp(local_pes_1_16_io_out_sum_exp),
    .io_out_kv(local_pes_1_16_io_out_kv),
    .io_out_stage(local_pes_1_16_io_out_stage)
  );
  PE_1 local_pes_1_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_17_clock),
    .reset(local_pes_1_17_reset),
    .io_in_q(local_pes_1_17_io_in_q),
    .io_in_sum(local_pes_1_17_io_in_sum),
    .io_in_sum_exp(local_pes_1_17_io_in_sum_exp),
    .io_in_kv(local_pes_1_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_17_io_in_inv_sum),
    .io_in_stage(local_pes_1_17_io_in_stage),
    .io_out_q(local_pes_1_17_io_out_q),
    .io_out_sum(local_pes_1_17_io_out_sum),
    .io_out_sum_exp(local_pes_1_17_io_out_sum_exp),
    .io_out_kv(local_pes_1_17_io_out_kv),
    .io_out_stage(local_pes_1_17_io_out_stage)
  );
  PE_1 local_pes_1_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_18_clock),
    .reset(local_pes_1_18_reset),
    .io_in_q(local_pes_1_18_io_in_q),
    .io_in_sum(local_pes_1_18_io_in_sum),
    .io_in_sum_exp(local_pes_1_18_io_in_sum_exp),
    .io_in_kv(local_pes_1_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_18_io_in_inv_sum),
    .io_in_stage(local_pes_1_18_io_in_stage),
    .io_out_q(local_pes_1_18_io_out_q),
    .io_out_sum(local_pes_1_18_io_out_sum),
    .io_out_sum_exp(local_pes_1_18_io_out_sum_exp),
    .io_out_kv(local_pes_1_18_io_out_kv),
    .io_out_stage(local_pes_1_18_io_out_stage)
  );
  PE_1 local_pes_1_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_19_clock),
    .reset(local_pes_1_19_reset),
    .io_in_q(local_pes_1_19_io_in_q),
    .io_in_sum(local_pes_1_19_io_in_sum),
    .io_in_sum_exp(local_pes_1_19_io_in_sum_exp),
    .io_in_kv(local_pes_1_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_19_io_in_inv_sum),
    .io_in_stage(local_pes_1_19_io_in_stage),
    .io_out_q(local_pes_1_19_io_out_q),
    .io_out_sum(local_pes_1_19_io_out_sum),
    .io_out_sum_exp(local_pes_1_19_io_out_sum_exp),
    .io_out_kv(local_pes_1_19_io_out_kv),
    .io_out_stage(local_pes_1_19_io_out_stage)
  );
  PE_1 local_pes_1_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_20_clock),
    .reset(local_pes_1_20_reset),
    .io_in_q(local_pes_1_20_io_in_q),
    .io_in_sum(local_pes_1_20_io_in_sum),
    .io_in_sum_exp(local_pes_1_20_io_in_sum_exp),
    .io_in_kv(local_pes_1_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_20_io_in_inv_sum),
    .io_in_stage(local_pes_1_20_io_in_stage),
    .io_out_q(local_pes_1_20_io_out_q),
    .io_out_sum(local_pes_1_20_io_out_sum),
    .io_out_sum_exp(local_pes_1_20_io_out_sum_exp),
    .io_out_kv(local_pes_1_20_io_out_kv),
    .io_out_stage(local_pes_1_20_io_out_stage)
  );
  PE_1 local_pes_1_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_21_clock),
    .reset(local_pes_1_21_reset),
    .io_in_q(local_pes_1_21_io_in_q),
    .io_in_sum(local_pes_1_21_io_in_sum),
    .io_in_sum_exp(local_pes_1_21_io_in_sum_exp),
    .io_in_kv(local_pes_1_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_21_io_in_inv_sum),
    .io_in_stage(local_pes_1_21_io_in_stage),
    .io_out_q(local_pes_1_21_io_out_q),
    .io_out_sum(local_pes_1_21_io_out_sum),
    .io_out_sum_exp(local_pes_1_21_io_out_sum_exp),
    .io_out_kv(local_pes_1_21_io_out_kv),
    .io_out_stage(local_pes_1_21_io_out_stage)
  );
  PE_1 local_pes_1_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_22_clock),
    .reset(local_pes_1_22_reset),
    .io_in_q(local_pes_1_22_io_in_q),
    .io_in_sum(local_pes_1_22_io_in_sum),
    .io_in_sum_exp(local_pes_1_22_io_in_sum_exp),
    .io_in_kv(local_pes_1_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_22_io_in_inv_sum),
    .io_in_stage(local_pes_1_22_io_in_stage),
    .io_out_q(local_pes_1_22_io_out_q),
    .io_out_sum(local_pes_1_22_io_out_sum),
    .io_out_sum_exp(local_pes_1_22_io_out_sum_exp),
    .io_out_kv(local_pes_1_22_io_out_kv),
    .io_out_stage(local_pes_1_22_io_out_stage)
  );
  PE_1 local_pes_1_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_23_clock),
    .reset(local_pes_1_23_reset),
    .io_in_q(local_pes_1_23_io_in_q),
    .io_in_sum(local_pes_1_23_io_in_sum),
    .io_in_sum_exp(local_pes_1_23_io_in_sum_exp),
    .io_in_kv(local_pes_1_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_23_io_in_inv_sum),
    .io_in_stage(local_pes_1_23_io_in_stage),
    .io_out_q(local_pes_1_23_io_out_q),
    .io_out_sum(local_pes_1_23_io_out_sum),
    .io_out_sum_exp(local_pes_1_23_io_out_sum_exp),
    .io_out_kv(local_pes_1_23_io_out_kv),
    .io_out_stage(local_pes_1_23_io_out_stage)
  );
  PE_1 local_pes_1_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_24_clock),
    .reset(local_pes_1_24_reset),
    .io_in_q(local_pes_1_24_io_in_q),
    .io_in_sum(local_pes_1_24_io_in_sum),
    .io_in_sum_exp(local_pes_1_24_io_in_sum_exp),
    .io_in_kv(local_pes_1_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_24_io_in_inv_sum),
    .io_in_stage(local_pes_1_24_io_in_stage),
    .io_out_q(local_pes_1_24_io_out_q),
    .io_out_sum(local_pes_1_24_io_out_sum),
    .io_out_sum_exp(local_pes_1_24_io_out_sum_exp),
    .io_out_kv(local_pes_1_24_io_out_kv),
    .io_out_stage(local_pes_1_24_io_out_stage)
  );
  PE_1 local_pes_1_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_25_clock),
    .reset(local_pes_1_25_reset),
    .io_in_q(local_pes_1_25_io_in_q),
    .io_in_sum(local_pes_1_25_io_in_sum),
    .io_in_sum_exp(local_pes_1_25_io_in_sum_exp),
    .io_in_kv(local_pes_1_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_25_io_in_inv_sum),
    .io_in_stage(local_pes_1_25_io_in_stage),
    .io_out_q(local_pes_1_25_io_out_q),
    .io_out_sum(local_pes_1_25_io_out_sum),
    .io_out_sum_exp(local_pes_1_25_io_out_sum_exp),
    .io_out_kv(local_pes_1_25_io_out_kv),
    .io_out_stage(local_pes_1_25_io_out_stage)
  );
  PE_1 local_pes_1_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_26_clock),
    .reset(local_pes_1_26_reset),
    .io_in_q(local_pes_1_26_io_in_q),
    .io_in_sum(local_pes_1_26_io_in_sum),
    .io_in_sum_exp(local_pes_1_26_io_in_sum_exp),
    .io_in_kv(local_pes_1_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_26_io_in_inv_sum),
    .io_in_stage(local_pes_1_26_io_in_stage),
    .io_out_q(local_pes_1_26_io_out_q),
    .io_out_sum(local_pes_1_26_io_out_sum),
    .io_out_sum_exp(local_pes_1_26_io_out_sum_exp),
    .io_out_kv(local_pes_1_26_io_out_kv),
    .io_out_stage(local_pes_1_26_io_out_stage)
  );
  PE_1 local_pes_1_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_27_clock),
    .reset(local_pes_1_27_reset),
    .io_in_q(local_pes_1_27_io_in_q),
    .io_in_sum(local_pes_1_27_io_in_sum),
    .io_in_sum_exp(local_pes_1_27_io_in_sum_exp),
    .io_in_kv(local_pes_1_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_27_io_in_inv_sum),
    .io_in_stage(local_pes_1_27_io_in_stage),
    .io_out_q(local_pes_1_27_io_out_q),
    .io_out_sum(local_pes_1_27_io_out_sum),
    .io_out_sum_exp(local_pes_1_27_io_out_sum_exp),
    .io_out_kv(local_pes_1_27_io_out_kv),
    .io_out_stage(local_pes_1_27_io_out_stage)
  );
  PE_1 local_pes_1_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_28_clock),
    .reset(local_pes_1_28_reset),
    .io_in_q(local_pes_1_28_io_in_q),
    .io_in_sum(local_pes_1_28_io_in_sum),
    .io_in_sum_exp(local_pes_1_28_io_in_sum_exp),
    .io_in_kv(local_pes_1_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_28_io_in_inv_sum),
    .io_in_stage(local_pes_1_28_io_in_stage),
    .io_out_q(local_pes_1_28_io_out_q),
    .io_out_sum(local_pes_1_28_io_out_sum),
    .io_out_sum_exp(local_pes_1_28_io_out_sum_exp),
    .io_out_kv(local_pes_1_28_io_out_kv),
    .io_out_stage(local_pes_1_28_io_out_stage)
  );
  PE_1 local_pes_1_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_29_clock),
    .reset(local_pes_1_29_reset),
    .io_in_q(local_pes_1_29_io_in_q),
    .io_in_sum(local_pes_1_29_io_in_sum),
    .io_in_sum_exp(local_pes_1_29_io_in_sum_exp),
    .io_in_kv(local_pes_1_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_29_io_in_inv_sum),
    .io_in_stage(local_pes_1_29_io_in_stage),
    .io_out_q(local_pes_1_29_io_out_q),
    .io_out_sum(local_pes_1_29_io_out_sum),
    .io_out_sum_exp(local_pes_1_29_io_out_sum_exp),
    .io_out_kv(local_pes_1_29_io_out_kv),
    .io_out_stage(local_pes_1_29_io_out_stage)
  );
  PE_1 local_pes_1_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_30_clock),
    .reset(local_pes_1_30_reset),
    .io_in_q(local_pes_1_30_io_in_q),
    .io_in_sum(local_pes_1_30_io_in_sum),
    .io_in_sum_exp(local_pes_1_30_io_in_sum_exp),
    .io_in_kv(local_pes_1_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_30_io_in_inv_sum),
    .io_in_stage(local_pes_1_30_io_in_stage),
    .io_out_q(local_pes_1_30_io_out_q),
    .io_out_sum(local_pes_1_30_io_out_sum),
    .io_out_sum_exp(local_pes_1_30_io_out_sum_exp),
    .io_out_kv(local_pes_1_30_io_out_kv),
    .io_out_stage(local_pes_1_30_io_out_stage)
  );
  PE_1 local_pes_1_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_1_31_clock),
    .reset(local_pes_1_31_reset),
    .io_in_q(local_pes_1_31_io_in_q),
    .io_in_sum(local_pes_1_31_io_in_sum),
    .io_in_sum_exp(local_pes_1_31_io_in_sum_exp),
    .io_in_kv(local_pes_1_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_1_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_1_31_io_in_inv_sum),
    .io_in_stage(local_pes_1_31_io_in_stage),
    .io_out_q(local_pes_1_31_io_out_q),
    .io_out_sum(local_pes_1_31_io_out_sum),
    .io_out_sum_exp(local_pes_1_31_io_out_sum_exp),
    .io_out_kv(local_pes_1_31_io_out_kv),
    .io_out_stage(local_pes_1_31_io_out_stage)
  );
  PE local_pes_2_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_0_clock),
    .reset(local_pes_2_0_reset),
    .io_in_q(local_pes_2_0_io_in_q),
    .io_in_kv(local_pes_2_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_0_io_in_inv_sum),
    .io_in_stage(local_pes_2_0_io_in_stage),
    .io_out_q(local_pes_2_0_io_out_q),
    .io_out_sum(local_pes_2_0_io_out_sum),
    .io_out_kv(local_pes_2_0_io_out_kv),
    .io_out_stage(local_pes_2_0_io_out_stage)
  );
  PE_1 local_pes_2_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_1_clock),
    .reset(local_pes_2_1_reset),
    .io_in_q(local_pes_2_1_io_in_q),
    .io_in_sum(local_pes_2_1_io_in_sum),
    .io_in_sum_exp(local_pes_2_1_io_in_sum_exp),
    .io_in_kv(local_pes_2_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_1_io_in_inv_sum),
    .io_in_stage(local_pes_2_1_io_in_stage),
    .io_out_q(local_pes_2_1_io_out_q),
    .io_out_sum(local_pes_2_1_io_out_sum),
    .io_out_sum_exp(local_pes_2_1_io_out_sum_exp),
    .io_out_kv(local_pes_2_1_io_out_kv),
    .io_out_stage(local_pes_2_1_io_out_stage)
  );
  PE_1 local_pes_2_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_2_clock),
    .reset(local_pes_2_2_reset),
    .io_in_q(local_pes_2_2_io_in_q),
    .io_in_sum(local_pes_2_2_io_in_sum),
    .io_in_sum_exp(local_pes_2_2_io_in_sum_exp),
    .io_in_kv(local_pes_2_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_2_io_in_inv_sum),
    .io_in_stage(local_pes_2_2_io_in_stage),
    .io_out_q(local_pes_2_2_io_out_q),
    .io_out_sum(local_pes_2_2_io_out_sum),
    .io_out_sum_exp(local_pes_2_2_io_out_sum_exp),
    .io_out_kv(local_pes_2_2_io_out_kv),
    .io_out_stage(local_pes_2_2_io_out_stage)
  );
  PE_1 local_pes_2_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_3_clock),
    .reset(local_pes_2_3_reset),
    .io_in_q(local_pes_2_3_io_in_q),
    .io_in_sum(local_pes_2_3_io_in_sum),
    .io_in_sum_exp(local_pes_2_3_io_in_sum_exp),
    .io_in_kv(local_pes_2_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_3_io_in_inv_sum),
    .io_in_stage(local_pes_2_3_io_in_stage),
    .io_out_q(local_pes_2_3_io_out_q),
    .io_out_sum(local_pes_2_3_io_out_sum),
    .io_out_sum_exp(local_pes_2_3_io_out_sum_exp),
    .io_out_kv(local_pes_2_3_io_out_kv),
    .io_out_stage(local_pes_2_3_io_out_stage)
  );
  PE_1 local_pes_2_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_4_clock),
    .reset(local_pes_2_4_reset),
    .io_in_q(local_pes_2_4_io_in_q),
    .io_in_sum(local_pes_2_4_io_in_sum),
    .io_in_sum_exp(local_pes_2_4_io_in_sum_exp),
    .io_in_kv(local_pes_2_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_4_io_in_inv_sum),
    .io_in_stage(local_pes_2_4_io_in_stage),
    .io_out_q(local_pes_2_4_io_out_q),
    .io_out_sum(local_pes_2_4_io_out_sum),
    .io_out_sum_exp(local_pes_2_4_io_out_sum_exp),
    .io_out_kv(local_pes_2_4_io_out_kv),
    .io_out_stage(local_pes_2_4_io_out_stage)
  );
  PE_1 local_pes_2_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_5_clock),
    .reset(local_pes_2_5_reset),
    .io_in_q(local_pes_2_5_io_in_q),
    .io_in_sum(local_pes_2_5_io_in_sum),
    .io_in_sum_exp(local_pes_2_5_io_in_sum_exp),
    .io_in_kv(local_pes_2_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_5_io_in_inv_sum),
    .io_in_stage(local_pes_2_5_io_in_stage),
    .io_out_q(local_pes_2_5_io_out_q),
    .io_out_sum(local_pes_2_5_io_out_sum),
    .io_out_sum_exp(local_pes_2_5_io_out_sum_exp),
    .io_out_kv(local_pes_2_5_io_out_kv),
    .io_out_stage(local_pes_2_5_io_out_stage)
  );
  PE_1 local_pes_2_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_6_clock),
    .reset(local_pes_2_6_reset),
    .io_in_q(local_pes_2_6_io_in_q),
    .io_in_sum(local_pes_2_6_io_in_sum),
    .io_in_sum_exp(local_pes_2_6_io_in_sum_exp),
    .io_in_kv(local_pes_2_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_6_io_in_inv_sum),
    .io_in_stage(local_pes_2_6_io_in_stage),
    .io_out_q(local_pes_2_6_io_out_q),
    .io_out_sum(local_pes_2_6_io_out_sum),
    .io_out_sum_exp(local_pes_2_6_io_out_sum_exp),
    .io_out_kv(local_pes_2_6_io_out_kv),
    .io_out_stage(local_pes_2_6_io_out_stage)
  );
  PE_1 local_pes_2_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_7_clock),
    .reset(local_pes_2_7_reset),
    .io_in_q(local_pes_2_7_io_in_q),
    .io_in_sum(local_pes_2_7_io_in_sum),
    .io_in_sum_exp(local_pes_2_7_io_in_sum_exp),
    .io_in_kv(local_pes_2_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_7_io_in_inv_sum),
    .io_in_stage(local_pes_2_7_io_in_stage),
    .io_out_q(local_pes_2_7_io_out_q),
    .io_out_sum(local_pes_2_7_io_out_sum),
    .io_out_sum_exp(local_pes_2_7_io_out_sum_exp),
    .io_out_kv(local_pes_2_7_io_out_kv),
    .io_out_stage(local_pes_2_7_io_out_stage)
  );
  PE_1 local_pes_2_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_8_clock),
    .reset(local_pes_2_8_reset),
    .io_in_q(local_pes_2_8_io_in_q),
    .io_in_sum(local_pes_2_8_io_in_sum),
    .io_in_sum_exp(local_pes_2_8_io_in_sum_exp),
    .io_in_kv(local_pes_2_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_8_io_in_inv_sum),
    .io_in_stage(local_pes_2_8_io_in_stage),
    .io_out_q(local_pes_2_8_io_out_q),
    .io_out_sum(local_pes_2_8_io_out_sum),
    .io_out_sum_exp(local_pes_2_8_io_out_sum_exp),
    .io_out_kv(local_pes_2_8_io_out_kv),
    .io_out_stage(local_pes_2_8_io_out_stage)
  );
  PE_1 local_pes_2_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_9_clock),
    .reset(local_pes_2_9_reset),
    .io_in_q(local_pes_2_9_io_in_q),
    .io_in_sum(local_pes_2_9_io_in_sum),
    .io_in_sum_exp(local_pes_2_9_io_in_sum_exp),
    .io_in_kv(local_pes_2_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_9_io_in_inv_sum),
    .io_in_stage(local_pes_2_9_io_in_stage),
    .io_out_q(local_pes_2_9_io_out_q),
    .io_out_sum(local_pes_2_9_io_out_sum),
    .io_out_sum_exp(local_pes_2_9_io_out_sum_exp),
    .io_out_kv(local_pes_2_9_io_out_kv),
    .io_out_stage(local_pes_2_9_io_out_stage)
  );
  PE_1 local_pes_2_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_10_clock),
    .reset(local_pes_2_10_reset),
    .io_in_q(local_pes_2_10_io_in_q),
    .io_in_sum(local_pes_2_10_io_in_sum),
    .io_in_sum_exp(local_pes_2_10_io_in_sum_exp),
    .io_in_kv(local_pes_2_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_10_io_in_inv_sum),
    .io_in_stage(local_pes_2_10_io_in_stage),
    .io_out_q(local_pes_2_10_io_out_q),
    .io_out_sum(local_pes_2_10_io_out_sum),
    .io_out_sum_exp(local_pes_2_10_io_out_sum_exp),
    .io_out_kv(local_pes_2_10_io_out_kv),
    .io_out_stage(local_pes_2_10_io_out_stage)
  );
  PE_1 local_pes_2_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_11_clock),
    .reset(local_pes_2_11_reset),
    .io_in_q(local_pes_2_11_io_in_q),
    .io_in_sum(local_pes_2_11_io_in_sum),
    .io_in_sum_exp(local_pes_2_11_io_in_sum_exp),
    .io_in_kv(local_pes_2_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_11_io_in_inv_sum),
    .io_in_stage(local_pes_2_11_io_in_stage),
    .io_out_q(local_pes_2_11_io_out_q),
    .io_out_sum(local_pes_2_11_io_out_sum),
    .io_out_sum_exp(local_pes_2_11_io_out_sum_exp),
    .io_out_kv(local_pes_2_11_io_out_kv),
    .io_out_stage(local_pes_2_11_io_out_stage)
  );
  PE_1 local_pes_2_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_12_clock),
    .reset(local_pes_2_12_reset),
    .io_in_q(local_pes_2_12_io_in_q),
    .io_in_sum(local_pes_2_12_io_in_sum),
    .io_in_sum_exp(local_pes_2_12_io_in_sum_exp),
    .io_in_kv(local_pes_2_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_12_io_in_inv_sum),
    .io_in_stage(local_pes_2_12_io_in_stage),
    .io_out_q(local_pes_2_12_io_out_q),
    .io_out_sum(local_pes_2_12_io_out_sum),
    .io_out_sum_exp(local_pes_2_12_io_out_sum_exp),
    .io_out_kv(local_pes_2_12_io_out_kv),
    .io_out_stage(local_pes_2_12_io_out_stage)
  );
  PE_1 local_pes_2_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_13_clock),
    .reset(local_pes_2_13_reset),
    .io_in_q(local_pes_2_13_io_in_q),
    .io_in_sum(local_pes_2_13_io_in_sum),
    .io_in_sum_exp(local_pes_2_13_io_in_sum_exp),
    .io_in_kv(local_pes_2_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_13_io_in_inv_sum),
    .io_in_stage(local_pes_2_13_io_in_stage),
    .io_out_q(local_pes_2_13_io_out_q),
    .io_out_sum(local_pes_2_13_io_out_sum),
    .io_out_sum_exp(local_pes_2_13_io_out_sum_exp),
    .io_out_kv(local_pes_2_13_io_out_kv),
    .io_out_stage(local_pes_2_13_io_out_stage)
  );
  PE_1 local_pes_2_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_14_clock),
    .reset(local_pes_2_14_reset),
    .io_in_q(local_pes_2_14_io_in_q),
    .io_in_sum(local_pes_2_14_io_in_sum),
    .io_in_sum_exp(local_pes_2_14_io_in_sum_exp),
    .io_in_kv(local_pes_2_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_14_io_in_inv_sum),
    .io_in_stage(local_pes_2_14_io_in_stage),
    .io_out_q(local_pes_2_14_io_out_q),
    .io_out_sum(local_pes_2_14_io_out_sum),
    .io_out_sum_exp(local_pes_2_14_io_out_sum_exp),
    .io_out_kv(local_pes_2_14_io_out_kv),
    .io_out_stage(local_pes_2_14_io_out_stage)
  );
  PE_1 local_pes_2_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_15_clock),
    .reset(local_pes_2_15_reset),
    .io_in_q(local_pes_2_15_io_in_q),
    .io_in_sum(local_pes_2_15_io_in_sum),
    .io_in_sum_exp(local_pes_2_15_io_in_sum_exp),
    .io_in_kv(local_pes_2_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_15_io_in_inv_sum),
    .io_in_stage(local_pes_2_15_io_in_stage),
    .io_out_q(local_pes_2_15_io_out_q),
    .io_out_sum(local_pes_2_15_io_out_sum),
    .io_out_sum_exp(local_pes_2_15_io_out_sum_exp),
    .io_out_kv(local_pes_2_15_io_out_kv),
    .io_out_stage(local_pes_2_15_io_out_stage)
  );
  PE_1 local_pes_2_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_16_clock),
    .reset(local_pes_2_16_reset),
    .io_in_q(local_pes_2_16_io_in_q),
    .io_in_sum(local_pes_2_16_io_in_sum),
    .io_in_sum_exp(local_pes_2_16_io_in_sum_exp),
    .io_in_kv(local_pes_2_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_16_io_in_inv_sum),
    .io_in_stage(local_pes_2_16_io_in_stage),
    .io_out_q(local_pes_2_16_io_out_q),
    .io_out_sum(local_pes_2_16_io_out_sum),
    .io_out_sum_exp(local_pes_2_16_io_out_sum_exp),
    .io_out_kv(local_pes_2_16_io_out_kv),
    .io_out_stage(local_pes_2_16_io_out_stage)
  );
  PE_1 local_pes_2_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_17_clock),
    .reset(local_pes_2_17_reset),
    .io_in_q(local_pes_2_17_io_in_q),
    .io_in_sum(local_pes_2_17_io_in_sum),
    .io_in_sum_exp(local_pes_2_17_io_in_sum_exp),
    .io_in_kv(local_pes_2_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_17_io_in_inv_sum),
    .io_in_stage(local_pes_2_17_io_in_stage),
    .io_out_q(local_pes_2_17_io_out_q),
    .io_out_sum(local_pes_2_17_io_out_sum),
    .io_out_sum_exp(local_pes_2_17_io_out_sum_exp),
    .io_out_kv(local_pes_2_17_io_out_kv),
    .io_out_stage(local_pes_2_17_io_out_stage)
  );
  PE_1 local_pes_2_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_18_clock),
    .reset(local_pes_2_18_reset),
    .io_in_q(local_pes_2_18_io_in_q),
    .io_in_sum(local_pes_2_18_io_in_sum),
    .io_in_sum_exp(local_pes_2_18_io_in_sum_exp),
    .io_in_kv(local_pes_2_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_18_io_in_inv_sum),
    .io_in_stage(local_pes_2_18_io_in_stage),
    .io_out_q(local_pes_2_18_io_out_q),
    .io_out_sum(local_pes_2_18_io_out_sum),
    .io_out_sum_exp(local_pes_2_18_io_out_sum_exp),
    .io_out_kv(local_pes_2_18_io_out_kv),
    .io_out_stage(local_pes_2_18_io_out_stage)
  );
  PE_1 local_pes_2_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_19_clock),
    .reset(local_pes_2_19_reset),
    .io_in_q(local_pes_2_19_io_in_q),
    .io_in_sum(local_pes_2_19_io_in_sum),
    .io_in_sum_exp(local_pes_2_19_io_in_sum_exp),
    .io_in_kv(local_pes_2_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_19_io_in_inv_sum),
    .io_in_stage(local_pes_2_19_io_in_stage),
    .io_out_q(local_pes_2_19_io_out_q),
    .io_out_sum(local_pes_2_19_io_out_sum),
    .io_out_sum_exp(local_pes_2_19_io_out_sum_exp),
    .io_out_kv(local_pes_2_19_io_out_kv),
    .io_out_stage(local_pes_2_19_io_out_stage)
  );
  PE_1 local_pes_2_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_20_clock),
    .reset(local_pes_2_20_reset),
    .io_in_q(local_pes_2_20_io_in_q),
    .io_in_sum(local_pes_2_20_io_in_sum),
    .io_in_sum_exp(local_pes_2_20_io_in_sum_exp),
    .io_in_kv(local_pes_2_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_20_io_in_inv_sum),
    .io_in_stage(local_pes_2_20_io_in_stage),
    .io_out_q(local_pes_2_20_io_out_q),
    .io_out_sum(local_pes_2_20_io_out_sum),
    .io_out_sum_exp(local_pes_2_20_io_out_sum_exp),
    .io_out_kv(local_pes_2_20_io_out_kv),
    .io_out_stage(local_pes_2_20_io_out_stage)
  );
  PE_1 local_pes_2_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_21_clock),
    .reset(local_pes_2_21_reset),
    .io_in_q(local_pes_2_21_io_in_q),
    .io_in_sum(local_pes_2_21_io_in_sum),
    .io_in_sum_exp(local_pes_2_21_io_in_sum_exp),
    .io_in_kv(local_pes_2_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_21_io_in_inv_sum),
    .io_in_stage(local_pes_2_21_io_in_stage),
    .io_out_q(local_pes_2_21_io_out_q),
    .io_out_sum(local_pes_2_21_io_out_sum),
    .io_out_sum_exp(local_pes_2_21_io_out_sum_exp),
    .io_out_kv(local_pes_2_21_io_out_kv),
    .io_out_stage(local_pes_2_21_io_out_stage)
  );
  PE_1 local_pes_2_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_22_clock),
    .reset(local_pes_2_22_reset),
    .io_in_q(local_pes_2_22_io_in_q),
    .io_in_sum(local_pes_2_22_io_in_sum),
    .io_in_sum_exp(local_pes_2_22_io_in_sum_exp),
    .io_in_kv(local_pes_2_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_22_io_in_inv_sum),
    .io_in_stage(local_pes_2_22_io_in_stage),
    .io_out_q(local_pes_2_22_io_out_q),
    .io_out_sum(local_pes_2_22_io_out_sum),
    .io_out_sum_exp(local_pes_2_22_io_out_sum_exp),
    .io_out_kv(local_pes_2_22_io_out_kv),
    .io_out_stage(local_pes_2_22_io_out_stage)
  );
  PE_1 local_pes_2_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_23_clock),
    .reset(local_pes_2_23_reset),
    .io_in_q(local_pes_2_23_io_in_q),
    .io_in_sum(local_pes_2_23_io_in_sum),
    .io_in_sum_exp(local_pes_2_23_io_in_sum_exp),
    .io_in_kv(local_pes_2_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_23_io_in_inv_sum),
    .io_in_stage(local_pes_2_23_io_in_stage),
    .io_out_q(local_pes_2_23_io_out_q),
    .io_out_sum(local_pes_2_23_io_out_sum),
    .io_out_sum_exp(local_pes_2_23_io_out_sum_exp),
    .io_out_kv(local_pes_2_23_io_out_kv),
    .io_out_stage(local_pes_2_23_io_out_stage)
  );
  PE_1 local_pes_2_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_24_clock),
    .reset(local_pes_2_24_reset),
    .io_in_q(local_pes_2_24_io_in_q),
    .io_in_sum(local_pes_2_24_io_in_sum),
    .io_in_sum_exp(local_pes_2_24_io_in_sum_exp),
    .io_in_kv(local_pes_2_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_24_io_in_inv_sum),
    .io_in_stage(local_pes_2_24_io_in_stage),
    .io_out_q(local_pes_2_24_io_out_q),
    .io_out_sum(local_pes_2_24_io_out_sum),
    .io_out_sum_exp(local_pes_2_24_io_out_sum_exp),
    .io_out_kv(local_pes_2_24_io_out_kv),
    .io_out_stage(local_pes_2_24_io_out_stage)
  );
  PE_1 local_pes_2_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_25_clock),
    .reset(local_pes_2_25_reset),
    .io_in_q(local_pes_2_25_io_in_q),
    .io_in_sum(local_pes_2_25_io_in_sum),
    .io_in_sum_exp(local_pes_2_25_io_in_sum_exp),
    .io_in_kv(local_pes_2_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_25_io_in_inv_sum),
    .io_in_stage(local_pes_2_25_io_in_stage),
    .io_out_q(local_pes_2_25_io_out_q),
    .io_out_sum(local_pes_2_25_io_out_sum),
    .io_out_sum_exp(local_pes_2_25_io_out_sum_exp),
    .io_out_kv(local_pes_2_25_io_out_kv),
    .io_out_stage(local_pes_2_25_io_out_stage)
  );
  PE_1 local_pes_2_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_26_clock),
    .reset(local_pes_2_26_reset),
    .io_in_q(local_pes_2_26_io_in_q),
    .io_in_sum(local_pes_2_26_io_in_sum),
    .io_in_sum_exp(local_pes_2_26_io_in_sum_exp),
    .io_in_kv(local_pes_2_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_26_io_in_inv_sum),
    .io_in_stage(local_pes_2_26_io_in_stage),
    .io_out_q(local_pes_2_26_io_out_q),
    .io_out_sum(local_pes_2_26_io_out_sum),
    .io_out_sum_exp(local_pes_2_26_io_out_sum_exp),
    .io_out_kv(local_pes_2_26_io_out_kv),
    .io_out_stage(local_pes_2_26_io_out_stage)
  );
  PE_1 local_pes_2_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_27_clock),
    .reset(local_pes_2_27_reset),
    .io_in_q(local_pes_2_27_io_in_q),
    .io_in_sum(local_pes_2_27_io_in_sum),
    .io_in_sum_exp(local_pes_2_27_io_in_sum_exp),
    .io_in_kv(local_pes_2_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_27_io_in_inv_sum),
    .io_in_stage(local_pes_2_27_io_in_stage),
    .io_out_q(local_pes_2_27_io_out_q),
    .io_out_sum(local_pes_2_27_io_out_sum),
    .io_out_sum_exp(local_pes_2_27_io_out_sum_exp),
    .io_out_kv(local_pes_2_27_io_out_kv),
    .io_out_stage(local_pes_2_27_io_out_stage)
  );
  PE_1 local_pes_2_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_28_clock),
    .reset(local_pes_2_28_reset),
    .io_in_q(local_pes_2_28_io_in_q),
    .io_in_sum(local_pes_2_28_io_in_sum),
    .io_in_sum_exp(local_pes_2_28_io_in_sum_exp),
    .io_in_kv(local_pes_2_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_28_io_in_inv_sum),
    .io_in_stage(local_pes_2_28_io_in_stage),
    .io_out_q(local_pes_2_28_io_out_q),
    .io_out_sum(local_pes_2_28_io_out_sum),
    .io_out_sum_exp(local_pes_2_28_io_out_sum_exp),
    .io_out_kv(local_pes_2_28_io_out_kv),
    .io_out_stage(local_pes_2_28_io_out_stage)
  );
  PE_1 local_pes_2_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_29_clock),
    .reset(local_pes_2_29_reset),
    .io_in_q(local_pes_2_29_io_in_q),
    .io_in_sum(local_pes_2_29_io_in_sum),
    .io_in_sum_exp(local_pes_2_29_io_in_sum_exp),
    .io_in_kv(local_pes_2_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_29_io_in_inv_sum),
    .io_in_stage(local_pes_2_29_io_in_stage),
    .io_out_q(local_pes_2_29_io_out_q),
    .io_out_sum(local_pes_2_29_io_out_sum),
    .io_out_sum_exp(local_pes_2_29_io_out_sum_exp),
    .io_out_kv(local_pes_2_29_io_out_kv),
    .io_out_stage(local_pes_2_29_io_out_stage)
  );
  PE_1 local_pes_2_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_30_clock),
    .reset(local_pes_2_30_reset),
    .io_in_q(local_pes_2_30_io_in_q),
    .io_in_sum(local_pes_2_30_io_in_sum),
    .io_in_sum_exp(local_pes_2_30_io_in_sum_exp),
    .io_in_kv(local_pes_2_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_30_io_in_inv_sum),
    .io_in_stage(local_pes_2_30_io_in_stage),
    .io_out_q(local_pes_2_30_io_out_q),
    .io_out_sum(local_pes_2_30_io_out_sum),
    .io_out_sum_exp(local_pes_2_30_io_out_sum_exp),
    .io_out_kv(local_pes_2_30_io_out_kv),
    .io_out_stage(local_pes_2_30_io_out_stage)
  );
  PE_1 local_pes_2_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_2_31_clock),
    .reset(local_pes_2_31_reset),
    .io_in_q(local_pes_2_31_io_in_q),
    .io_in_sum(local_pes_2_31_io_in_sum),
    .io_in_sum_exp(local_pes_2_31_io_in_sum_exp),
    .io_in_kv(local_pes_2_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_2_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_2_31_io_in_inv_sum),
    .io_in_stage(local_pes_2_31_io_in_stage),
    .io_out_q(local_pes_2_31_io_out_q),
    .io_out_sum(local_pes_2_31_io_out_sum),
    .io_out_sum_exp(local_pes_2_31_io_out_sum_exp),
    .io_out_kv(local_pes_2_31_io_out_kv),
    .io_out_stage(local_pes_2_31_io_out_stage)
  );
  PE local_pes_3_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_0_clock),
    .reset(local_pes_3_0_reset),
    .io_in_q(local_pes_3_0_io_in_q),
    .io_in_kv(local_pes_3_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_0_io_in_inv_sum),
    .io_in_stage(local_pes_3_0_io_in_stage),
    .io_out_q(local_pes_3_0_io_out_q),
    .io_out_sum(local_pes_3_0_io_out_sum),
    .io_out_kv(local_pes_3_0_io_out_kv),
    .io_out_stage(local_pes_3_0_io_out_stage)
  );
  PE_1 local_pes_3_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_1_clock),
    .reset(local_pes_3_1_reset),
    .io_in_q(local_pes_3_1_io_in_q),
    .io_in_sum(local_pes_3_1_io_in_sum),
    .io_in_sum_exp(local_pes_3_1_io_in_sum_exp),
    .io_in_kv(local_pes_3_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_1_io_in_inv_sum),
    .io_in_stage(local_pes_3_1_io_in_stage),
    .io_out_q(local_pes_3_1_io_out_q),
    .io_out_sum(local_pes_3_1_io_out_sum),
    .io_out_sum_exp(local_pes_3_1_io_out_sum_exp),
    .io_out_kv(local_pes_3_1_io_out_kv),
    .io_out_stage(local_pes_3_1_io_out_stage)
  );
  PE_1 local_pes_3_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_2_clock),
    .reset(local_pes_3_2_reset),
    .io_in_q(local_pes_3_2_io_in_q),
    .io_in_sum(local_pes_3_2_io_in_sum),
    .io_in_sum_exp(local_pes_3_2_io_in_sum_exp),
    .io_in_kv(local_pes_3_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_2_io_in_inv_sum),
    .io_in_stage(local_pes_3_2_io_in_stage),
    .io_out_q(local_pes_3_2_io_out_q),
    .io_out_sum(local_pes_3_2_io_out_sum),
    .io_out_sum_exp(local_pes_3_2_io_out_sum_exp),
    .io_out_kv(local_pes_3_2_io_out_kv),
    .io_out_stage(local_pes_3_2_io_out_stage)
  );
  PE_1 local_pes_3_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_3_clock),
    .reset(local_pes_3_3_reset),
    .io_in_q(local_pes_3_3_io_in_q),
    .io_in_sum(local_pes_3_3_io_in_sum),
    .io_in_sum_exp(local_pes_3_3_io_in_sum_exp),
    .io_in_kv(local_pes_3_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_3_io_in_inv_sum),
    .io_in_stage(local_pes_3_3_io_in_stage),
    .io_out_q(local_pes_3_3_io_out_q),
    .io_out_sum(local_pes_3_3_io_out_sum),
    .io_out_sum_exp(local_pes_3_3_io_out_sum_exp),
    .io_out_kv(local_pes_3_3_io_out_kv),
    .io_out_stage(local_pes_3_3_io_out_stage)
  );
  PE_1 local_pes_3_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_4_clock),
    .reset(local_pes_3_4_reset),
    .io_in_q(local_pes_3_4_io_in_q),
    .io_in_sum(local_pes_3_4_io_in_sum),
    .io_in_sum_exp(local_pes_3_4_io_in_sum_exp),
    .io_in_kv(local_pes_3_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_4_io_in_inv_sum),
    .io_in_stage(local_pes_3_4_io_in_stage),
    .io_out_q(local_pes_3_4_io_out_q),
    .io_out_sum(local_pes_3_4_io_out_sum),
    .io_out_sum_exp(local_pes_3_4_io_out_sum_exp),
    .io_out_kv(local_pes_3_4_io_out_kv),
    .io_out_stage(local_pes_3_4_io_out_stage)
  );
  PE_1 local_pes_3_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_5_clock),
    .reset(local_pes_3_5_reset),
    .io_in_q(local_pes_3_5_io_in_q),
    .io_in_sum(local_pes_3_5_io_in_sum),
    .io_in_sum_exp(local_pes_3_5_io_in_sum_exp),
    .io_in_kv(local_pes_3_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_5_io_in_inv_sum),
    .io_in_stage(local_pes_3_5_io_in_stage),
    .io_out_q(local_pes_3_5_io_out_q),
    .io_out_sum(local_pes_3_5_io_out_sum),
    .io_out_sum_exp(local_pes_3_5_io_out_sum_exp),
    .io_out_kv(local_pes_3_5_io_out_kv),
    .io_out_stage(local_pes_3_5_io_out_stage)
  );
  PE_1 local_pes_3_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_6_clock),
    .reset(local_pes_3_6_reset),
    .io_in_q(local_pes_3_6_io_in_q),
    .io_in_sum(local_pes_3_6_io_in_sum),
    .io_in_sum_exp(local_pes_3_6_io_in_sum_exp),
    .io_in_kv(local_pes_3_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_6_io_in_inv_sum),
    .io_in_stage(local_pes_3_6_io_in_stage),
    .io_out_q(local_pes_3_6_io_out_q),
    .io_out_sum(local_pes_3_6_io_out_sum),
    .io_out_sum_exp(local_pes_3_6_io_out_sum_exp),
    .io_out_kv(local_pes_3_6_io_out_kv),
    .io_out_stage(local_pes_3_6_io_out_stage)
  );
  PE_1 local_pes_3_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_7_clock),
    .reset(local_pes_3_7_reset),
    .io_in_q(local_pes_3_7_io_in_q),
    .io_in_sum(local_pes_3_7_io_in_sum),
    .io_in_sum_exp(local_pes_3_7_io_in_sum_exp),
    .io_in_kv(local_pes_3_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_7_io_in_inv_sum),
    .io_in_stage(local_pes_3_7_io_in_stage),
    .io_out_q(local_pes_3_7_io_out_q),
    .io_out_sum(local_pes_3_7_io_out_sum),
    .io_out_sum_exp(local_pes_3_7_io_out_sum_exp),
    .io_out_kv(local_pes_3_7_io_out_kv),
    .io_out_stage(local_pes_3_7_io_out_stage)
  );
  PE_1 local_pes_3_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_8_clock),
    .reset(local_pes_3_8_reset),
    .io_in_q(local_pes_3_8_io_in_q),
    .io_in_sum(local_pes_3_8_io_in_sum),
    .io_in_sum_exp(local_pes_3_8_io_in_sum_exp),
    .io_in_kv(local_pes_3_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_8_io_in_inv_sum),
    .io_in_stage(local_pes_3_8_io_in_stage),
    .io_out_q(local_pes_3_8_io_out_q),
    .io_out_sum(local_pes_3_8_io_out_sum),
    .io_out_sum_exp(local_pes_3_8_io_out_sum_exp),
    .io_out_kv(local_pes_3_8_io_out_kv),
    .io_out_stage(local_pes_3_8_io_out_stage)
  );
  PE_1 local_pes_3_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_9_clock),
    .reset(local_pes_3_9_reset),
    .io_in_q(local_pes_3_9_io_in_q),
    .io_in_sum(local_pes_3_9_io_in_sum),
    .io_in_sum_exp(local_pes_3_9_io_in_sum_exp),
    .io_in_kv(local_pes_3_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_9_io_in_inv_sum),
    .io_in_stage(local_pes_3_9_io_in_stage),
    .io_out_q(local_pes_3_9_io_out_q),
    .io_out_sum(local_pes_3_9_io_out_sum),
    .io_out_sum_exp(local_pes_3_9_io_out_sum_exp),
    .io_out_kv(local_pes_3_9_io_out_kv),
    .io_out_stage(local_pes_3_9_io_out_stage)
  );
  PE_1 local_pes_3_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_10_clock),
    .reset(local_pes_3_10_reset),
    .io_in_q(local_pes_3_10_io_in_q),
    .io_in_sum(local_pes_3_10_io_in_sum),
    .io_in_sum_exp(local_pes_3_10_io_in_sum_exp),
    .io_in_kv(local_pes_3_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_10_io_in_inv_sum),
    .io_in_stage(local_pes_3_10_io_in_stage),
    .io_out_q(local_pes_3_10_io_out_q),
    .io_out_sum(local_pes_3_10_io_out_sum),
    .io_out_sum_exp(local_pes_3_10_io_out_sum_exp),
    .io_out_kv(local_pes_3_10_io_out_kv),
    .io_out_stage(local_pes_3_10_io_out_stage)
  );
  PE_1 local_pes_3_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_11_clock),
    .reset(local_pes_3_11_reset),
    .io_in_q(local_pes_3_11_io_in_q),
    .io_in_sum(local_pes_3_11_io_in_sum),
    .io_in_sum_exp(local_pes_3_11_io_in_sum_exp),
    .io_in_kv(local_pes_3_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_11_io_in_inv_sum),
    .io_in_stage(local_pes_3_11_io_in_stage),
    .io_out_q(local_pes_3_11_io_out_q),
    .io_out_sum(local_pes_3_11_io_out_sum),
    .io_out_sum_exp(local_pes_3_11_io_out_sum_exp),
    .io_out_kv(local_pes_3_11_io_out_kv),
    .io_out_stage(local_pes_3_11_io_out_stage)
  );
  PE_1 local_pes_3_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_12_clock),
    .reset(local_pes_3_12_reset),
    .io_in_q(local_pes_3_12_io_in_q),
    .io_in_sum(local_pes_3_12_io_in_sum),
    .io_in_sum_exp(local_pes_3_12_io_in_sum_exp),
    .io_in_kv(local_pes_3_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_12_io_in_inv_sum),
    .io_in_stage(local_pes_3_12_io_in_stage),
    .io_out_q(local_pes_3_12_io_out_q),
    .io_out_sum(local_pes_3_12_io_out_sum),
    .io_out_sum_exp(local_pes_3_12_io_out_sum_exp),
    .io_out_kv(local_pes_3_12_io_out_kv),
    .io_out_stage(local_pes_3_12_io_out_stage)
  );
  PE_1 local_pes_3_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_13_clock),
    .reset(local_pes_3_13_reset),
    .io_in_q(local_pes_3_13_io_in_q),
    .io_in_sum(local_pes_3_13_io_in_sum),
    .io_in_sum_exp(local_pes_3_13_io_in_sum_exp),
    .io_in_kv(local_pes_3_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_13_io_in_inv_sum),
    .io_in_stage(local_pes_3_13_io_in_stage),
    .io_out_q(local_pes_3_13_io_out_q),
    .io_out_sum(local_pes_3_13_io_out_sum),
    .io_out_sum_exp(local_pes_3_13_io_out_sum_exp),
    .io_out_kv(local_pes_3_13_io_out_kv),
    .io_out_stage(local_pes_3_13_io_out_stage)
  );
  PE_1 local_pes_3_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_14_clock),
    .reset(local_pes_3_14_reset),
    .io_in_q(local_pes_3_14_io_in_q),
    .io_in_sum(local_pes_3_14_io_in_sum),
    .io_in_sum_exp(local_pes_3_14_io_in_sum_exp),
    .io_in_kv(local_pes_3_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_14_io_in_inv_sum),
    .io_in_stage(local_pes_3_14_io_in_stage),
    .io_out_q(local_pes_3_14_io_out_q),
    .io_out_sum(local_pes_3_14_io_out_sum),
    .io_out_sum_exp(local_pes_3_14_io_out_sum_exp),
    .io_out_kv(local_pes_3_14_io_out_kv),
    .io_out_stage(local_pes_3_14_io_out_stage)
  );
  PE_1 local_pes_3_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_15_clock),
    .reset(local_pes_3_15_reset),
    .io_in_q(local_pes_3_15_io_in_q),
    .io_in_sum(local_pes_3_15_io_in_sum),
    .io_in_sum_exp(local_pes_3_15_io_in_sum_exp),
    .io_in_kv(local_pes_3_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_15_io_in_inv_sum),
    .io_in_stage(local_pes_3_15_io_in_stage),
    .io_out_q(local_pes_3_15_io_out_q),
    .io_out_sum(local_pes_3_15_io_out_sum),
    .io_out_sum_exp(local_pes_3_15_io_out_sum_exp),
    .io_out_kv(local_pes_3_15_io_out_kv),
    .io_out_stage(local_pes_3_15_io_out_stage)
  );
  PE_1 local_pes_3_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_16_clock),
    .reset(local_pes_3_16_reset),
    .io_in_q(local_pes_3_16_io_in_q),
    .io_in_sum(local_pes_3_16_io_in_sum),
    .io_in_sum_exp(local_pes_3_16_io_in_sum_exp),
    .io_in_kv(local_pes_3_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_16_io_in_inv_sum),
    .io_in_stage(local_pes_3_16_io_in_stage),
    .io_out_q(local_pes_3_16_io_out_q),
    .io_out_sum(local_pes_3_16_io_out_sum),
    .io_out_sum_exp(local_pes_3_16_io_out_sum_exp),
    .io_out_kv(local_pes_3_16_io_out_kv),
    .io_out_stage(local_pes_3_16_io_out_stage)
  );
  PE_1 local_pes_3_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_17_clock),
    .reset(local_pes_3_17_reset),
    .io_in_q(local_pes_3_17_io_in_q),
    .io_in_sum(local_pes_3_17_io_in_sum),
    .io_in_sum_exp(local_pes_3_17_io_in_sum_exp),
    .io_in_kv(local_pes_3_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_17_io_in_inv_sum),
    .io_in_stage(local_pes_3_17_io_in_stage),
    .io_out_q(local_pes_3_17_io_out_q),
    .io_out_sum(local_pes_3_17_io_out_sum),
    .io_out_sum_exp(local_pes_3_17_io_out_sum_exp),
    .io_out_kv(local_pes_3_17_io_out_kv),
    .io_out_stage(local_pes_3_17_io_out_stage)
  );
  PE_1 local_pes_3_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_18_clock),
    .reset(local_pes_3_18_reset),
    .io_in_q(local_pes_3_18_io_in_q),
    .io_in_sum(local_pes_3_18_io_in_sum),
    .io_in_sum_exp(local_pes_3_18_io_in_sum_exp),
    .io_in_kv(local_pes_3_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_18_io_in_inv_sum),
    .io_in_stage(local_pes_3_18_io_in_stage),
    .io_out_q(local_pes_3_18_io_out_q),
    .io_out_sum(local_pes_3_18_io_out_sum),
    .io_out_sum_exp(local_pes_3_18_io_out_sum_exp),
    .io_out_kv(local_pes_3_18_io_out_kv),
    .io_out_stage(local_pes_3_18_io_out_stage)
  );
  PE_1 local_pes_3_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_19_clock),
    .reset(local_pes_3_19_reset),
    .io_in_q(local_pes_3_19_io_in_q),
    .io_in_sum(local_pes_3_19_io_in_sum),
    .io_in_sum_exp(local_pes_3_19_io_in_sum_exp),
    .io_in_kv(local_pes_3_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_19_io_in_inv_sum),
    .io_in_stage(local_pes_3_19_io_in_stage),
    .io_out_q(local_pes_3_19_io_out_q),
    .io_out_sum(local_pes_3_19_io_out_sum),
    .io_out_sum_exp(local_pes_3_19_io_out_sum_exp),
    .io_out_kv(local_pes_3_19_io_out_kv),
    .io_out_stage(local_pes_3_19_io_out_stage)
  );
  PE_1 local_pes_3_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_20_clock),
    .reset(local_pes_3_20_reset),
    .io_in_q(local_pes_3_20_io_in_q),
    .io_in_sum(local_pes_3_20_io_in_sum),
    .io_in_sum_exp(local_pes_3_20_io_in_sum_exp),
    .io_in_kv(local_pes_3_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_20_io_in_inv_sum),
    .io_in_stage(local_pes_3_20_io_in_stage),
    .io_out_q(local_pes_3_20_io_out_q),
    .io_out_sum(local_pes_3_20_io_out_sum),
    .io_out_sum_exp(local_pes_3_20_io_out_sum_exp),
    .io_out_kv(local_pes_3_20_io_out_kv),
    .io_out_stage(local_pes_3_20_io_out_stage)
  );
  PE_1 local_pes_3_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_21_clock),
    .reset(local_pes_3_21_reset),
    .io_in_q(local_pes_3_21_io_in_q),
    .io_in_sum(local_pes_3_21_io_in_sum),
    .io_in_sum_exp(local_pes_3_21_io_in_sum_exp),
    .io_in_kv(local_pes_3_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_21_io_in_inv_sum),
    .io_in_stage(local_pes_3_21_io_in_stage),
    .io_out_q(local_pes_3_21_io_out_q),
    .io_out_sum(local_pes_3_21_io_out_sum),
    .io_out_sum_exp(local_pes_3_21_io_out_sum_exp),
    .io_out_kv(local_pes_3_21_io_out_kv),
    .io_out_stage(local_pes_3_21_io_out_stage)
  );
  PE_1 local_pes_3_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_22_clock),
    .reset(local_pes_3_22_reset),
    .io_in_q(local_pes_3_22_io_in_q),
    .io_in_sum(local_pes_3_22_io_in_sum),
    .io_in_sum_exp(local_pes_3_22_io_in_sum_exp),
    .io_in_kv(local_pes_3_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_22_io_in_inv_sum),
    .io_in_stage(local_pes_3_22_io_in_stage),
    .io_out_q(local_pes_3_22_io_out_q),
    .io_out_sum(local_pes_3_22_io_out_sum),
    .io_out_sum_exp(local_pes_3_22_io_out_sum_exp),
    .io_out_kv(local_pes_3_22_io_out_kv),
    .io_out_stage(local_pes_3_22_io_out_stage)
  );
  PE_1 local_pes_3_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_23_clock),
    .reset(local_pes_3_23_reset),
    .io_in_q(local_pes_3_23_io_in_q),
    .io_in_sum(local_pes_3_23_io_in_sum),
    .io_in_sum_exp(local_pes_3_23_io_in_sum_exp),
    .io_in_kv(local_pes_3_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_23_io_in_inv_sum),
    .io_in_stage(local_pes_3_23_io_in_stage),
    .io_out_q(local_pes_3_23_io_out_q),
    .io_out_sum(local_pes_3_23_io_out_sum),
    .io_out_sum_exp(local_pes_3_23_io_out_sum_exp),
    .io_out_kv(local_pes_3_23_io_out_kv),
    .io_out_stage(local_pes_3_23_io_out_stage)
  );
  PE_1 local_pes_3_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_24_clock),
    .reset(local_pes_3_24_reset),
    .io_in_q(local_pes_3_24_io_in_q),
    .io_in_sum(local_pes_3_24_io_in_sum),
    .io_in_sum_exp(local_pes_3_24_io_in_sum_exp),
    .io_in_kv(local_pes_3_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_24_io_in_inv_sum),
    .io_in_stage(local_pes_3_24_io_in_stage),
    .io_out_q(local_pes_3_24_io_out_q),
    .io_out_sum(local_pes_3_24_io_out_sum),
    .io_out_sum_exp(local_pes_3_24_io_out_sum_exp),
    .io_out_kv(local_pes_3_24_io_out_kv),
    .io_out_stage(local_pes_3_24_io_out_stage)
  );
  PE_1 local_pes_3_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_25_clock),
    .reset(local_pes_3_25_reset),
    .io_in_q(local_pes_3_25_io_in_q),
    .io_in_sum(local_pes_3_25_io_in_sum),
    .io_in_sum_exp(local_pes_3_25_io_in_sum_exp),
    .io_in_kv(local_pes_3_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_25_io_in_inv_sum),
    .io_in_stage(local_pes_3_25_io_in_stage),
    .io_out_q(local_pes_3_25_io_out_q),
    .io_out_sum(local_pes_3_25_io_out_sum),
    .io_out_sum_exp(local_pes_3_25_io_out_sum_exp),
    .io_out_kv(local_pes_3_25_io_out_kv),
    .io_out_stage(local_pes_3_25_io_out_stage)
  );
  PE_1 local_pes_3_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_26_clock),
    .reset(local_pes_3_26_reset),
    .io_in_q(local_pes_3_26_io_in_q),
    .io_in_sum(local_pes_3_26_io_in_sum),
    .io_in_sum_exp(local_pes_3_26_io_in_sum_exp),
    .io_in_kv(local_pes_3_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_26_io_in_inv_sum),
    .io_in_stage(local_pes_3_26_io_in_stage),
    .io_out_q(local_pes_3_26_io_out_q),
    .io_out_sum(local_pes_3_26_io_out_sum),
    .io_out_sum_exp(local_pes_3_26_io_out_sum_exp),
    .io_out_kv(local_pes_3_26_io_out_kv),
    .io_out_stage(local_pes_3_26_io_out_stage)
  );
  PE_1 local_pes_3_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_27_clock),
    .reset(local_pes_3_27_reset),
    .io_in_q(local_pes_3_27_io_in_q),
    .io_in_sum(local_pes_3_27_io_in_sum),
    .io_in_sum_exp(local_pes_3_27_io_in_sum_exp),
    .io_in_kv(local_pes_3_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_27_io_in_inv_sum),
    .io_in_stage(local_pes_3_27_io_in_stage),
    .io_out_q(local_pes_3_27_io_out_q),
    .io_out_sum(local_pes_3_27_io_out_sum),
    .io_out_sum_exp(local_pes_3_27_io_out_sum_exp),
    .io_out_kv(local_pes_3_27_io_out_kv),
    .io_out_stage(local_pes_3_27_io_out_stage)
  );
  PE_1 local_pes_3_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_28_clock),
    .reset(local_pes_3_28_reset),
    .io_in_q(local_pes_3_28_io_in_q),
    .io_in_sum(local_pes_3_28_io_in_sum),
    .io_in_sum_exp(local_pes_3_28_io_in_sum_exp),
    .io_in_kv(local_pes_3_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_28_io_in_inv_sum),
    .io_in_stage(local_pes_3_28_io_in_stage),
    .io_out_q(local_pes_3_28_io_out_q),
    .io_out_sum(local_pes_3_28_io_out_sum),
    .io_out_sum_exp(local_pes_3_28_io_out_sum_exp),
    .io_out_kv(local_pes_3_28_io_out_kv),
    .io_out_stage(local_pes_3_28_io_out_stage)
  );
  PE_1 local_pes_3_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_29_clock),
    .reset(local_pes_3_29_reset),
    .io_in_q(local_pes_3_29_io_in_q),
    .io_in_sum(local_pes_3_29_io_in_sum),
    .io_in_sum_exp(local_pes_3_29_io_in_sum_exp),
    .io_in_kv(local_pes_3_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_29_io_in_inv_sum),
    .io_in_stage(local_pes_3_29_io_in_stage),
    .io_out_q(local_pes_3_29_io_out_q),
    .io_out_sum(local_pes_3_29_io_out_sum),
    .io_out_sum_exp(local_pes_3_29_io_out_sum_exp),
    .io_out_kv(local_pes_3_29_io_out_kv),
    .io_out_stage(local_pes_3_29_io_out_stage)
  );
  PE_1 local_pes_3_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_30_clock),
    .reset(local_pes_3_30_reset),
    .io_in_q(local_pes_3_30_io_in_q),
    .io_in_sum(local_pes_3_30_io_in_sum),
    .io_in_sum_exp(local_pes_3_30_io_in_sum_exp),
    .io_in_kv(local_pes_3_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_30_io_in_inv_sum),
    .io_in_stage(local_pes_3_30_io_in_stage),
    .io_out_q(local_pes_3_30_io_out_q),
    .io_out_sum(local_pes_3_30_io_out_sum),
    .io_out_sum_exp(local_pes_3_30_io_out_sum_exp),
    .io_out_kv(local_pes_3_30_io_out_kv),
    .io_out_stage(local_pes_3_30_io_out_stage)
  );
  PE_1 local_pes_3_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_3_31_clock),
    .reset(local_pes_3_31_reset),
    .io_in_q(local_pes_3_31_io_in_q),
    .io_in_sum(local_pes_3_31_io_in_sum),
    .io_in_sum_exp(local_pes_3_31_io_in_sum_exp),
    .io_in_kv(local_pes_3_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_3_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_3_31_io_in_inv_sum),
    .io_in_stage(local_pes_3_31_io_in_stage),
    .io_out_q(local_pes_3_31_io_out_q),
    .io_out_sum(local_pes_3_31_io_out_sum),
    .io_out_sum_exp(local_pes_3_31_io_out_sum_exp),
    .io_out_kv(local_pes_3_31_io_out_kv),
    .io_out_stage(local_pes_3_31_io_out_stage)
  );
  PE local_pes_4_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_0_clock),
    .reset(local_pes_4_0_reset),
    .io_in_q(local_pes_4_0_io_in_q),
    .io_in_kv(local_pes_4_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_0_io_in_inv_sum),
    .io_in_stage(local_pes_4_0_io_in_stage),
    .io_out_q(local_pes_4_0_io_out_q),
    .io_out_sum(local_pes_4_0_io_out_sum),
    .io_out_kv(local_pes_4_0_io_out_kv),
    .io_out_stage(local_pes_4_0_io_out_stage)
  );
  PE_1 local_pes_4_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_1_clock),
    .reset(local_pes_4_1_reset),
    .io_in_q(local_pes_4_1_io_in_q),
    .io_in_sum(local_pes_4_1_io_in_sum),
    .io_in_sum_exp(local_pes_4_1_io_in_sum_exp),
    .io_in_kv(local_pes_4_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_1_io_in_inv_sum),
    .io_in_stage(local_pes_4_1_io_in_stage),
    .io_out_q(local_pes_4_1_io_out_q),
    .io_out_sum(local_pes_4_1_io_out_sum),
    .io_out_sum_exp(local_pes_4_1_io_out_sum_exp),
    .io_out_kv(local_pes_4_1_io_out_kv),
    .io_out_stage(local_pes_4_1_io_out_stage)
  );
  PE_1 local_pes_4_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_2_clock),
    .reset(local_pes_4_2_reset),
    .io_in_q(local_pes_4_2_io_in_q),
    .io_in_sum(local_pes_4_2_io_in_sum),
    .io_in_sum_exp(local_pes_4_2_io_in_sum_exp),
    .io_in_kv(local_pes_4_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_2_io_in_inv_sum),
    .io_in_stage(local_pes_4_2_io_in_stage),
    .io_out_q(local_pes_4_2_io_out_q),
    .io_out_sum(local_pes_4_2_io_out_sum),
    .io_out_sum_exp(local_pes_4_2_io_out_sum_exp),
    .io_out_kv(local_pes_4_2_io_out_kv),
    .io_out_stage(local_pes_4_2_io_out_stage)
  );
  PE_1 local_pes_4_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_3_clock),
    .reset(local_pes_4_3_reset),
    .io_in_q(local_pes_4_3_io_in_q),
    .io_in_sum(local_pes_4_3_io_in_sum),
    .io_in_sum_exp(local_pes_4_3_io_in_sum_exp),
    .io_in_kv(local_pes_4_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_3_io_in_inv_sum),
    .io_in_stage(local_pes_4_3_io_in_stage),
    .io_out_q(local_pes_4_3_io_out_q),
    .io_out_sum(local_pes_4_3_io_out_sum),
    .io_out_sum_exp(local_pes_4_3_io_out_sum_exp),
    .io_out_kv(local_pes_4_3_io_out_kv),
    .io_out_stage(local_pes_4_3_io_out_stage)
  );
  PE_1 local_pes_4_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_4_clock),
    .reset(local_pes_4_4_reset),
    .io_in_q(local_pes_4_4_io_in_q),
    .io_in_sum(local_pes_4_4_io_in_sum),
    .io_in_sum_exp(local_pes_4_4_io_in_sum_exp),
    .io_in_kv(local_pes_4_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_4_io_in_inv_sum),
    .io_in_stage(local_pes_4_4_io_in_stage),
    .io_out_q(local_pes_4_4_io_out_q),
    .io_out_sum(local_pes_4_4_io_out_sum),
    .io_out_sum_exp(local_pes_4_4_io_out_sum_exp),
    .io_out_kv(local_pes_4_4_io_out_kv),
    .io_out_stage(local_pes_4_4_io_out_stage)
  );
  PE_1 local_pes_4_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_5_clock),
    .reset(local_pes_4_5_reset),
    .io_in_q(local_pes_4_5_io_in_q),
    .io_in_sum(local_pes_4_5_io_in_sum),
    .io_in_sum_exp(local_pes_4_5_io_in_sum_exp),
    .io_in_kv(local_pes_4_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_5_io_in_inv_sum),
    .io_in_stage(local_pes_4_5_io_in_stage),
    .io_out_q(local_pes_4_5_io_out_q),
    .io_out_sum(local_pes_4_5_io_out_sum),
    .io_out_sum_exp(local_pes_4_5_io_out_sum_exp),
    .io_out_kv(local_pes_4_5_io_out_kv),
    .io_out_stage(local_pes_4_5_io_out_stage)
  );
  PE_1 local_pes_4_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_6_clock),
    .reset(local_pes_4_6_reset),
    .io_in_q(local_pes_4_6_io_in_q),
    .io_in_sum(local_pes_4_6_io_in_sum),
    .io_in_sum_exp(local_pes_4_6_io_in_sum_exp),
    .io_in_kv(local_pes_4_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_6_io_in_inv_sum),
    .io_in_stage(local_pes_4_6_io_in_stage),
    .io_out_q(local_pes_4_6_io_out_q),
    .io_out_sum(local_pes_4_6_io_out_sum),
    .io_out_sum_exp(local_pes_4_6_io_out_sum_exp),
    .io_out_kv(local_pes_4_6_io_out_kv),
    .io_out_stage(local_pes_4_6_io_out_stage)
  );
  PE_1 local_pes_4_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_7_clock),
    .reset(local_pes_4_7_reset),
    .io_in_q(local_pes_4_7_io_in_q),
    .io_in_sum(local_pes_4_7_io_in_sum),
    .io_in_sum_exp(local_pes_4_7_io_in_sum_exp),
    .io_in_kv(local_pes_4_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_7_io_in_inv_sum),
    .io_in_stage(local_pes_4_7_io_in_stage),
    .io_out_q(local_pes_4_7_io_out_q),
    .io_out_sum(local_pes_4_7_io_out_sum),
    .io_out_sum_exp(local_pes_4_7_io_out_sum_exp),
    .io_out_kv(local_pes_4_7_io_out_kv),
    .io_out_stage(local_pes_4_7_io_out_stage)
  );
  PE_1 local_pes_4_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_8_clock),
    .reset(local_pes_4_8_reset),
    .io_in_q(local_pes_4_8_io_in_q),
    .io_in_sum(local_pes_4_8_io_in_sum),
    .io_in_sum_exp(local_pes_4_8_io_in_sum_exp),
    .io_in_kv(local_pes_4_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_8_io_in_inv_sum),
    .io_in_stage(local_pes_4_8_io_in_stage),
    .io_out_q(local_pes_4_8_io_out_q),
    .io_out_sum(local_pes_4_8_io_out_sum),
    .io_out_sum_exp(local_pes_4_8_io_out_sum_exp),
    .io_out_kv(local_pes_4_8_io_out_kv),
    .io_out_stage(local_pes_4_8_io_out_stage)
  );
  PE_1 local_pes_4_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_9_clock),
    .reset(local_pes_4_9_reset),
    .io_in_q(local_pes_4_9_io_in_q),
    .io_in_sum(local_pes_4_9_io_in_sum),
    .io_in_sum_exp(local_pes_4_9_io_in_sum_exp),
    .io_in_kv(local_pes_4_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_9_io_in_inv_sum),
    .io_in_stage(local_pes_4_9_io_in_stage),
    .io_out_q(local_pes_4_9_io_out_q),
    .io_out_sum(local_pes_4_9_io_out_sum),
    .io_out_sum_exp(local_pes_4_9_io_out_sum_exp),
    .io_out_kv(local_pes_4_9_io_out_kv),
    .io_out_stage(local_pes_4_9_io_out_stage)
  );
  PE_1 local_pes_4_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_10_clock),
    .reset(local_pes_4_10_reset),
    .io_in_q(local_pes_4_10_io_in_q),
    .io_in_sum(local_pes_4_10_io_in_sum),
    .io_in_sum_exp(local_pes_4_10_io_in_sum_exp),
    .io_in_kv(local_pes_4_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_10_io_in_inv_sum),
    .io_in_stage(local_pes_4_10_io_in_stage),
    .io_out_q(local_pes_4_10_io_out_q),
    .io_out_sum(local_pes_4_10_io_out_sum),
    .io_out_sum_exp(local_pes_4_10_io_out_sum_exp),
    .io_out_kv(local_pes_4_10_io_out_kv),
    .io_out_stage(local_pes_4_10_io_out_stage)
  );
  PE_1 local_pes_4_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_11_clock),
    .reset(local_pes_4_11_reset),
    .io_in_q(local_pes_4_11_io_in_q),
    .io_in_sum(local_pes_4_11_io_in_sum),
    .io_in_sum_exp(local_pes_4_11_io_in_sum_exp),
    .io_in_kv(local_pes_4_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_11_io_in_inv_sum),
    .io_in_stage(local_pes_4_11_io_in_stage),
    .io_out_q(local_pes_4_11_io_out_q),
    .io_out_sum(local_pes_4_11_io_out_sum),
    .io_out_sum_exp(local_pes_4_11_io_out_sum_exp),
    .io_out_kv(local_pes_4_11_io_out_kv),
    .io_out_stage(local_pes_4_11_io_out_stage)
  );
  PE_1 local_pes_4_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_12_clock),
    .reset(local_pes_4_12_reset),
    .io_in_q(local_pes_4_12_io_in_q),
    .io_in_sum(local_pes_4_12_io_in_sum),
    .io_in_sum_exp(local_pes_4_12_io_in_sum_exp),
    .io_in_kv(local_pes_4_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_12_io_in_inv_sum),
    .io_in_stage(local_pes_4_12_io_in_stage),
    .io_out_q(local_pes_4_12_io_out_q),
    .io_out_sum(local_pes_4_12_io_out_sum),
    .io_out_sum_exp(local_pes_4_12_io_out_sum_exp),
    .io_out_kv(local_pes_4_12_io_out_kv),
    .io_out_stage(local_pes_4_12_io_out_stage)
  );
  PE_1 local_pes_4_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_13_clock),
    .reset(local_pes_4_13_reset),
    .io_in_q(local_pes_4_13_io_in_q),
    .io_in_sum(local_pes_4_13_io_in_sum),
    .io_in_sum_exp(local_pes_4_13_io_in_sum_exp),
    .io_in_kv(local_pes_4_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_13_io_in_inv_sum),
    .io_in_stage(local_pes_4_13_io_in_stage),
    .io_out_q(local_pes_4_13_io_out_q),
    .io_out_sum(local_pes_4_13_io_out_sum),
    .io_out_sum_exp(local_pes_4_13_io_out_sum_exp),
    .io_out_kv(local_pes_4_13_io_out_kv),
    .io_out_stage(local_pes_4_13_io_out_stage)
  );
  PE_1 local_pes_4_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_14_clock),
    .reset(local_pes_4_14_reset),
    .io_in_q(local_pes_4_14_io_in_q),
    .io_in_sum(local_pes_4_14_io_in_sum),
    .io_in_sum_exp(local_pes_4_14_io_in_sum_exp),
    .io_in_kv(local_pes_4_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_14_io_in_inv_sum),
    .io_in_stage(local_pes_4_14_io_in_stage),
    .io_out_q(local_pes_4_14_io_out_q),
    .io_out_sum(local_pes_4_14_io_out_sum),
    .io_out_sum_exp(local_pes_4_14_io_out_sum_exp),
    .io_out_kv(local_pes_4_14_io_out_kv),
    .io_out_stage(local_pes_4_14_io_out_stage)
  );
  PE_1 local_pes_4_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_15_clock),
    .reset(local_pes_4_15_reset),
    .io_in_q(local_pes_4_15_io_in_q),
    .io_in_sum(local_pes_4_15_io_in_sum),
    .io_in_sum_exp(local_pes_4_15_io_in_sum_exp),
    .io_in_kv(local_pes_4_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_15_io_in_inv_sum),
    .io_in_stage(local_pes_4_15_io_in_stage),
    .io_out_q(local_pes_4_15_io_out_q),
    .io_out_sum(local_pes_4_15_io_out_sum),
    .io_out_sum_exp(local_pes_4_15_io_out_sum_exp),
    .io_out_kv(local_pes_4_15_io_out_kv),
    .io_out_stage(local_pes_4_15_io_out_stage)
  );
  PE_1 local_pes_4_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_16_clock),
    .reset(local_pes_4_16_reset),
    .io_in_q(local_pes_4_16_io_in_q),
    .io_in_sum(local_pes_4_16_io_in_sum),
    .io_in_sum_exp(local_pes_4_16_io_in_sum_exp),
    .io_in_kv(local_pes_4_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_16_io_in_inv_sum),
    .io_in_stage(local_pes_4_16_io_in_stage),
    .io_out_q(local_pes_4_16_io_out_q),
    .io_out_sum(local_pes_4_16_io_out_sum),
    .io_out_sum_exp(local_pes_4_16_io_out_sum_exp),
    .io_out_kv(local_pes_4_16_io_out_kv),
    .io_out_stage(local_pes_4_16_io_out_stage)
  );
  PE_1 local_pes_4_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_17_clock),
    .reset(local_pes_4_17_reset),
    .io_in_q(local_pes_4_17_io_in_q),
    .io_in_sum(local_pes_4_17_io_in_sum),
    .io_in_sum_exp(local_pes_4_17_io_in_sum_exp),
    .io_in_kv(local_pes_4_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_17_io_in_inv_sum),
    .io_in_stage(local_pes_4_17_io_in_stage),
    .io_out_q(local_pes_4_17_io_out_q),
    .io_out_sum(local_pes_4_17_io_out_sum),
    .io_out_sum_exp(local_pes_4_17_io_out_sum_exp),
    .io_out_kv(local_pes_4_17_io_out_kv),
    .io_out_stage(local_pes_4_17_io_out_stage)
  );
  PE_1 local_pes_4_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_18_clock),
    .reset(local_pes_4_18_reset),
    .io_in_q(local_pes_4_18_io_in_q),
    .io_in_sum(local_pes_4_18_io_in_sum),
    .io_in_sum_exp(local_pes_4_18_io_in_sum_exp),
    .io_in_kv(local_pes_4_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_18_io_in_inv_sum),
    .io_in_stage(local_pes_4_18_io_in_stage),
    .io_out_q(local_pes_4_18_io_out_q),
    .io_out_sum(local_pes_4_18_io_out_sum),
    .io_out_sum_exp(local_pes_4_18_io_out_sum_exp),
    .io_out_kv(local_pes_4_18_io_out_kv),
    .io_out_stage(local_pes_4_18_io_out_stage)
  );
  PE_1 local_pes_4_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_19_clock),
    .reset(local_pes_4_19_reset),
    .io_in_q(local_pes_4_19_io_in_q),
    .io_in_sum(local_pes_4_19_io_in_sum),
    .io_in_sum_exp(local_pes_4_19_io_in_sum_exp),
    .io_in_kv(local_pes_4_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_19_io_in_inv_sum),
    .io_in_stage(local_pes_4_19_io_in_stage),
    .io_out_q(local_pes_4_19_io_out_q),
    .io_out_sum(local_pes_4_19_io_out_sum),
    .io_out_sum_exp(local_pes_4_19_io_out_sum_exp),
    .io_out_kv(local_pes_4_19_io_out_kv),
    .io_out_stage(local_pes_4_19_io_out_stage)
  );
  PE_1 local_pes_4_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_20_clock),
    .reset(local_pes_4_20_reset),
    .io_in_q(local_pes_4_20_io_in_q),
    .io_in_sum(local_pes_4_20_io_in_sum),
    .io_in_sum_exp(local_pes_4_20_io_in_sum_exp),
    .io_in_kv(local_pes_4_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_20_io_in_inv_sum),
    .io_in_stage(local_pes_4_20_io_in_stage),
    .io_out_q(local_pes_4_20_io_out_q),
    .io_out_sum(local_pes_4_20_io_out_sum),
    .io_out_sum_exp(local_pes_4_20_io_out_sum_exp),
    .io_out_kv(local_pes_4_20_io_out_kv),
    .io_out_stage(local_pes_4_20_io_out_stage)
  );
  PE_1 local_pes_4_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_21_clock),
    .reset(local_pes_4_21_reset),
    .io_in_q(local_pes_4_21_io_in_q),
    .io_in_sum(local_pes_4_21_io_in_sum),
    .io_in_sum_exp(local_pes_4_21_io_in_sum_exp),
    .io_in_kv(local_pes_4_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_21_io_in_inv_sum),
    .io_in_stage(local_pes_4_21_io_in_stage),
    .io_out_q(local_pes_4_21_io_out_q),
    .io_out_sum(local_pes_4_21_io_out_sum),
    .io_out_sum_exp(local_pes_4_21_io_out_sum_exp),
    .io_out_kv(local_pes_4_21_io_out_kv),
    .io_out_stage(local_pes_4_21_io_out_stage)
  );
  PE_1 local_pes_4_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_22_clock),
    .reset(local_pes_4_22_reset),
    .io_in_q(local_pes_4_22_io_in_q),
    .io_in_sum(local_pes_4_22_io_in_sum),
    .io_in_sum_exp(local_pes_4_22_io_in_sum_exp),
    .io_in_kv(local_pes_4_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_22_io_in_inv_sum),
    .io_in_stage(local_pes_4_22_io_in_stage),
    .io_out_q(local_pes_4_22_io_out_q),
    .io_out_sum(local_pes_4_22_io_out_sum),
    .io_out_sum_exp(local_pes_4_22_io_out_sum_exp),
    .io_out_kv(local_pes_4_22_io_out_kv),
    .io_out_stage(local_pes_4_22_io_out_stage)
  );
  PE_1 local_pes_4_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_23_clock),
    .reset(local_pes_4_23_reset),
    .io_in_q(local_pes_4_23_io_in_q),
    .io_in_sum(local_pes_4_23_io_in_sum),
    .io_in_sum_exp(local_pes_4_23_io_in_sum_exp),
    .io_in_kv(local_pes_4_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_23_io_in_inv_sum),
    .io_in_stage(local_pes_4_23_io_in_stage),
    .io_out_q(local_pes_4_23_io_out_q),
    .io_out_sum(local_pes_4_23_io_out_sum),
    .io_out_sum_exp(local_pes_4_23_io_out_sum_exp),
    .io_out_kv(local_pes_4_23_io_out_kv),
    .io_out_stage(local_pes_4_23_io_out_stage)
  );
  PE_1 local_pes_4_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_24_clock),
    .reset(local_pes_4_24_reset),
    .io_in_q(local_pes_4_24_io_in_q),
    .io_in_sum(local_pes_4_24_io_in_sum),
    .io_in_sum_exp(local_pes_4_24_io_in_sum_exp),
    .io_in_kv(local_pes_4_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_24_io_in_inv_sum),
    .io_in_stage(local_pes_4_24_io_in_stage),
    .io_out_q(local_pes_4_24_io_out_q),
    .io_out_sum(local_pes_4_24_io_out_sum),
    .io_out_sum_exp(local_pes_4_24_io_out_sum_exp),
    .io_out_kv(local_pes_4_24_io_out_kv),
    .io_out_stage(local_pes_4_24_io_out_stage)
  );
  PE_1 local_pes_4_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_25_clock),
    .reset(local_pes_4_25_reset),
    .io_in_q(local_pes_4_25_io_in_q),
    .io_in_sum(local_pes_4_25_io_in_sum),
    .io_in_sum_exp(local_pes_4_25_io_in_sum_exp),
    .io_in_kv(local_pes_4_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_25_io_in_inv_sum),
    .io_in_stage(local_pes_4_25_io_in_stage),
    .io_out_q(local_pes_4_25_io_out_q),
    .io_out_sum(local_pes_4_25_io_out_sum),
    .io_out_sum_exp(local_pes_4_25_io_out_sum_exp),
    .io_out_kv(local_pes_4_25_io_out_kv),
    .io_out_stage(local_pes_4_25_io_out_stage)
  );
  PE_1 local_pes_4_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_26_clock),
    .reset(local_pes_4_26_reset),
    .io_in_q(local_pes_4_26_io_in_q),
    .io_in_sum(local_pes_4_26_io_in_sum),
    .io_in_sum_exp(local_pes_4_26_io_in_sum_exp),
    .io_in_kv(local_pes_4_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_26_io_in_inv_sum),
    .io_in_stage(local_pes_4_26_io_in_stage),
    .io_out_q(local_pes_4_26_io_out_q),
    .io_out_sum(local_pes_4_26_io_out_sum),
    .io_out_sum_exp(local_pes_4_26_io_out_sum_exp),
    .io_out_kv(local_pes_4_26_io_out_kv),
    .io_out_stage(local_pes_4_26_io_out_stage)
  );
  PE_1 local_pes_4_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_27_clock),
    .reset(local_pes_4_27_reset),
    .io_in_q(local_pes_4_27_io_in_q),
    .io_in_sum(local_pes_4_27_io_in_sum),
    .io_in_sum_exp(local_pes_4_27_io_in_sum_exp),
    .io_in_kv(local_pes_4_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_27_io_in_inv_sum),
    .io_in_stage(local_pes_4_27_io_in_stage),
    .io_out_q(local_pes_4_27_io_out_q),
    .io_out_sum(local_pes_4_27_io_out_sum),
    .io_out_sum_exp(local_pes_4_27_io_out_sum_exp),
    .io_out_kv(local_pes_4_27_io_out_kv),
    .io_out_stage(local_pes_4_27_io_out_stage)
  );
  PE_1 local_pes_4_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_28_clock),
    .reset(local_pes_4_28_reset),
    .io_in_q(local_pes_4_28_io_in_q),
    .io_in_sum(local_pes_4_28_io_in_sum),
    .io_in_sum_exp(local_pes_4_28_io_in_sum_exp),
    .io_in_kv(local_pes_4_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_28_io_in_inv_sum),
    .io_in_stage(local_pes_4_28_io_in_stage),
    .io_out_q(local_pes_4_28_io_out_q),
    .io_out_sum(local_pes_4_28_io_out_sum),
    .io_out_sum_exp(local_pes_4_28_io_out_sum_exp),
    .io_out_kv(local_pes_4_28_io_out_kv),
    .io_out_stage(local_pes_4_28_io_out_stage)
  );
  PE_1 local_pes_4_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_29_clock),
    .reset(local_pes_4_29_reset),
    .io_in_q(local_pes_4_29_io_in_q),
    .io_in_sum(local_pes_4_29_io_in_sum),
    .io_in_sum_exp(local_pes_4_29_io_in_sum_exp),
    .io_in_kv(local_pes_4_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_29_io_in_inv_sum),
    .io_in_stage(local_pes_4_29_io_in_stage),
    .io_out_q(local_pes_4_29_io_out_q),
    .io_out_sum(local_pes_4_29_io_out_sum),
    .io_out_sum_exp(local_pes_4_29_io_out_sum_exp),
    .io_out_kv(local_pes_4_29_io_out_kv),
    .io_out_stage(local_pes_4_29_io_out_stage)
  );
  PE_1 local_pes_4_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_30_clock),
    .reset(local_pes_4_30_reset),
    .io_in_q(local_pes_4_30_io_in_q),
    .io_in_sum(local_pes_4_30_io_in_sum),
    .io_in_sum_exp(local_pes_4_30_io_in_sum_exp),
    .io_in_kv(local_pes_4_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_30_io_in_inv_sum),
    .io_in_stage(local_pes_4_30_io_in_stage),
    .io_out_q(local_pes_4_30_io_out_q),
    .io_out_sum(local_pes_4_30_io_out_sum),
    .io_out_sum_exp(local_pes_4_30_io_out_sum_exp),
    .io_out_kv(local_pes_4_30_io_out_kv),
    .io_out_stage(local_pes_4_30_io_out_stage)
  );
  PE_1 local_pes_4_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_4_31_clock),
    .reset(local_pes_4_31_reset),
    .io_in_q(local_pes_4_31_io_in_q),
    .io_in_sum(local_pes_4_31_io_in_sum),
    .io_in_sum_exp(local_pes_4_31_io_in_sum_exp),
    .io_in_kv(local_pes_4_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_4_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_4_31_io_in_inv_sum),
    .io_in_stage(local_pes_4_31_io_in_stage),
    .io_out_q(local_pes_4_31_io_out_q),
    .io_out_sum(local_pes_4_31_io_out_sum),
    .io_out_sum_exp(local_pes_4_31_io_out_sum_exp),
    .io_out_kv(local_pes_4_31_io_out_kv),
    .io_out_stage(local_pes_4_31_io_out_stage)
  );
  PE local_pes_5_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_0_clock),
    .reset(local_pes_5_0_reset),
    .io_in_q(local_pes_5_0_io_in_q),
    .io_in_kv(local_pes_5_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_0_io_in_inv_sum),
    .io_in_stage(local_pes_5_0_io_in_stage),
    .io_out_q(local_pes_5_0_io_out_q),
    .io_out_sum(local_pes_5_0_io_out_sum),
    .io_out_kv(local_pes_5_0_io_out_kv),
    .io_out_stage(local_pes_5_0_io_out_stage)
  );
  PE_1 local_pes_5_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_1_clock),
    .reset(local_pes_5_1_reset),
    .io_in_q(local_pes_5_1_io_in_q),
    .io_in_sum(local_pes_5_1_io_in_sum),
    .io_in_sum_exp(local_pes_5_1_io_in_sum_exp),
    .io_in_kv(local_pes_5_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_1_io_in_inv_sum),
    .io_in_stage(local_pes_5_1_io_in_stage),
    .io_out_q(local_pes_5_1_io_out_q),
    .io_out_sum(local_pes_5_1_io_out_sum),
    .io_out_sum_exp(local_pes_5_1_io_out_sum_exp),
    .io_out_kv(local_pes_5_1_io_out_kv),
    .io_out_stage(local_pes_5_1_io_out_stage)
  );
  PE_1 local_pes_5_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_2_clock),
    .reset(local_pes_5_2_reset),
    .io_in_q(local_pes_5_2_io_in_q),
    .io_in_sum(local_pes_5_2_io_in_sum),
    .io_in_sum_exp(local_pes_5_2_io_in_sum_exp),
    .io_in_kv(local_pes_5_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_2_io_in_inv_sum),
    .io_in_stage(local_pes_5_2_io_in_stage),
    .io_out_q(local_pes_5_2_io_out_q),
    .io_out_sum(local_pes_5_2_io_out_sum),
    .io_out_sum_exp(local_pes_5_2_io_out_sum_exp),
    .io_out_kv(local_pes_5_2_io_out_kv),
    .io_out_stage(local_pes_5_2_io_out_stage)
  );
  PE_1 local_pes_5_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_3_clock),
    .reset(local_pes_5_3_reset),
    .io_in_q(local_pes_5_3_io_in_q),
    .io_in_sum(local_pes_5_3_io_in_sum),
    .io_in_sum_exp(local_pes_5_3_io_in_sum_exp),
    .io_in_kv(local_pes_5_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_3_io_in_inv_sum),
    .io_in_stage(local_pes_5_3_io_in_stage),
    .io_out_q(local_pes_5_3_io_out_q),
    .io_out_sum(local_pes_5_3_io_out_sum),
    .io_out_sum_exp(local_pes_5_3_io_out_sum_exp),
    .io_out_kv(local_pes_5_3_io_out_kv),
    .io_out_stage(local_pes_5_3_io_out_stage)
  );
  PE_1 local_pes_5_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_4_clock),
    .reset(local_pes_5_4_reset),
    .io_in_q(local_pes_5_4_io_in_q),
    .io_in_sum(local_pes_5_4_io_in_sum),
    .io_in_sum_exp(local_pes_5_4_io_in_sum_exp),
    .io_in_kv(local_pes_5_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_4_io_in_inv_sum),
    .io_in_stage(local_pes_5_4_io_in_stage),
    .io_out_q(local_pes_5_4_io_out_q),
    .io_out_sum(local_pes_5_4_io_out_sum),
    .io_out_sum_exp(local_pes_5_4_io_out_sum_exp),
    .io_out_kv(local_pes_5_4_io_out_kv),
    .io_out_stage(local_pes_5_4_io_out_stage)
  );
  PE_1 local_pes_5_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_5_clock),
    .reset(local_pes_5_5_reset),
    .io_in_q(local_pes_5_5_io_in_q),
    .io_in_sum(local_pes_5_5_io_in_sum),
    .io_in_sum_exp(local_pes_5_5_io_in_sum_exp),
    .io_in_kv(local_pes_5_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_5_io_in_inv_sum),
    .io_in_stage(local_pes_5_5_io_in_stage),
    .io_out_q(local_pes_5_5_io_out_q),
    .io_out_sum(local_pes_5_5_io_out_sum),
    .io_out_sum_exp(local_pes_5_5_io_out_sum_exp),
    .io_out_kv(local_pes_5_5_io_out_kv),
    .io_out_stage(local_pes_5_5_io_out_stage)
  );
  PE_1 local_pes_5_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_6_clock),
    .reset(local_pes_5_6_reset),
    .io_in_q(local_pes_5_6_io_in_q),
    .io_in_sum(local_pes_5_6_io_in_sum),
    .io_in_sum_exp(local_pes_5_6_io_in_sum_exp),
    .io_in_kv(local_pes_5_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_6_io_in_inv_sum),
    .io_in_stage(local_pes_5_6_io_in_stage),
    .io_out_q(local_pes_5_6_io_out_q),
    .io_out_sum(local_pes_5_6_io_out_sum),
    .io_out_sum_exp(local_pes_5_6_io_out_sum_exp),
    .io_out_kv(local_pes_5_6_io_out_kv),
    .io_out_stage(local_pes_5_6_io_out_stage)
  );
  PE_1 local_pes_5_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_7_clock),
    .reset(local_pes_5_7_reset),
    .io_in_q(local_pes_5_7_io_in_q),
    .io_in_sum(local_pes_5_7_io_in_sum),
    .io_in_sum_exp(local_pes_5_7_io_in_sum_exp),
    .io_in_kv(local_pes_5_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_7_io_in_inv_sum),
    .io_in_stage(local_pes_5_7_io_in_stage),
    .io_out_q(local_pes_5_7_io_out_q),
    .io_out_sum(local_pes_5_7_io_out_sum),
    .io_out_sum_exp(local_pes_5_7_io_out_sum_exp),
    .io_out_kv(local_pes_5_7_io_out_kv),
    .io_out_stage(local_pes_5_7_io_out_stage)
  );
  PE_1 local_pes_5_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_8_clock),
    .reset(local_pes_5_8_reset),
    .io_in_q(local_pes_5_8_io_in_q),
    .io_in_sum(local_pes_5_8_io_in_sum),
    .io_in_sum_exp(local_pes_5_8_io_in_sum_exp),
    .io_in_kv(local_pes_5_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_8_io_in_inv_sum),
    .io_in_stage(local_pes_5_8_io_in_stage),
    .io_out_q(local_pes_5_8_io_out_q),
    .io_out_sum(local_pes_5_8_io_out_sum),
    .io_out_sum_exp(local_pes_5_8_io_out_sum_exp),
    .io_out_kv(local_pes_5_8_io_out_kv),
    .io_out_stage(local_pes_5_8_io_out_stage)
  );
  PE_1 local_pes_5_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_9_clock),
    .reset(local_pes_5_9_reset),
    .io_in_q(local_pes_5_9_io_in_q),
    .io_in_sum(local_pes_5_9_io_in_sum),
    .io_in_sum_exp(local_pes_5_9_io_in_sum_exp),
    .io_in_kv(local_pes_5_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_9_io_in_inv_sum),
    .io_in_stage(local_pes_5_9_io_in_stage),
    .io_out_q(local_pes_5_9_io_out_q),
    .io_out_sum(local_pes_5_9_io_out_sum),
    .io_out_sum_exp(local_pes_5_9_io_out_sum_exp),
    .io_out_kv(local_pes_5_9_io_out_kv),
    .io_out_stage(local_pes_5_9_io_out_stage)
  );
  PE_1 local_pes_5_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_10_clock),
    .reset(local_pes_5_10_reset),
    .io_in_q(local_pes_5_10_io_in_q),
    .io_in_sum(local_pes_5_10_io_in_sum),
    .io_in_sum_exp(local_pes_5_10_io_in_sum_exp),
    .io_in_kv(local_pes_5_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_10_io_in_inv_sum),
    .io_in_stage(local_pes_5_10_io_in_stage),
    .io_out_q(local_pes_5_10_io_out_q),
    .io_out_sum(local_pes_5_10_io_out_sum),
    .io_out_sum_exp(local_pes_5_10_io_out_sum_exp),
    .io_out_kv(local_pes_5_10_io_out_kv),
    .io_out_stage(local_pes_5_10_io_out_stage)
  );
  PE_1 local_pes_5_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_11_clock),
    .reset(local_pes_5_11_reset),
    .io_in_q(local_pes_5_11_io_in_q),
    .io_in_sum(local_pes_5_11_io_in_sum),
    .io_in_sum_exp(local_pes_5_11_io_in_sum_exp),
    .io_in_kv(local_pes_5_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_11_io_in_inv_sum),
    .io_in_stage(local_pes_5_11_io_in_stage),
    .io_out_q(local_pes_5_11_io_out_q),
    .io_out_sum(local_pes_5_11_io_out_sum),
    .io_out_sum_exp(local_pes_5_11_io_out_sum_exp),
    .io_out_kv(local_pes_5_11_io_out_kv),
    .io_out_stage(local_pes_5_11_io_out_stage)
  );
  PE_1 local_pes_5_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_12_clock),
    .reset(local_pes_5_12_reset),
    .io_in_q(local_pes_5_12_io_in_q),
    .io_in_sum(local_pes_5_12_io_in_sum),
    .io_in_sum_exp(local_pes_5_12_io_in_sum_exp),
    .io_in_kv(local_pes_5_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_12_io_in_inv_sum),
    .io_in_stage(local_pes_5_12_io_in_stage),
    .io_out_q(local_pes_5_12_io_out_q),
    .io_out_sum(local_pes_5_12_io_out_sum),
    .io_out_sum_exp(local_pes_5_12_io_out_sum_exp),
    .io_out_kv(local_pes_5_12_io_out_kv),
    .io_out_stage(local_pes_5_12_io_out_stage)
  );
  PE_1 local_pes_5_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_13_clock),
    .reset(local_pes_5_13_reset),
    .io_in_q(local_pes_5_13_io_in_q),
    .io_in_sum(local_pes_5_13_io_in_sum),
    .io_in_sum_exp(local_pes_5_13_io_in_sum_exp),
    .io_in_kv(local_pes_5_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_13_io_in_inv_sum),
    .io_in_stage(local_pes_5_13_io_in_stage),
    .io_out_q(local_pes_5_13_io_out_q),
    .io_out_sum(local_pes_5_13_io_out_sum),
    .io_out_sum_exp(local_pes_5_13_io_out_sum_exp),
    .io_out_kv(local_pes_5_13_io_out_kv),
    .io_out_stage(local_pes_5_13_io_out_stage)
  );
  PE_1 local_pes_5_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_14_clock),
    .reset(local_pes_5_14_reset),
    .io_in_q(local_pes_5_14_io_in_q),
    .io_in_sum(local_pes_5_14_io_in_sum),
    .io_in_sum_exp(local_pes_5_14_io_in_sum_exp),
    .io_in_kv(local_pes_5_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_14_io_in_inv_sum),
    .io_in_stage(local_pes_5_14_io_in_stage),
    .io_out_q(local_pes_5_14_io_out_q),
    .io_out_sum(local_pes_5_14_io_out_sum),
    .io_out_sum_exp(local_pes_5_14_io_out_sum_exp),
    .io_out_kv(local_pes_5_14_io_out_kv),
    .io_out_stage(local_pes_5_14_io_out_stage)
  );
  PE_1 local_pes_5_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_15_clock),
    .reset(local_pes_5_15_reset),
    .io_in_q(local_pes_5_15_io_in_q),
    .io_in_sum(local_pes_5_15_io_in_sum),
    .io_in_sum_exp(local_pes_5_15_io_in_sum_exp),
    .io_in_kv(local_pes_5_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_15_io_in_inv_sum),
    .io_in_stage(local_pes_5_15_io_in_stage),
    .io_out_q(local_pes_5_15_io_out_q),
    .io_out_sum(local_pes_5_15_io_out_sum),
    .io_out_sum_exp(local_pes_5_15_io_out_sum_exp),
    .io_out_kv(local_pes_5_15_io_out_kv),
    .io_out_stage(local_pes_5_15_io_out_stage)
  );
  PE_1 local_pes_5_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_16_clock),
    .reset(local_pes_5_16_reset),
    .io_in_q(local_pes_5_16_io_in_q),
    .io_in_sum(local_pes_5_16_io_in_sum),
    .io_in_sum_exp(local_pes_5_16_io_in_sum_exp),
    .io_in_kv(local_pes_5_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_16_io_in_inv_sum),
    .io_in_stage(local_pes_5_16_io_in_stage),
    .io_out_q(local_pes_5_16_io_out_q),
    .io_out_sum(local_pes_5_16_io_out_sum),
    .io_out_sum_exp(local_pes_5_16_io_out_sum_exp),
    .io_out_kv(local_pes_5_16_io_out_kv),
    .io_out_stage(local_pes_5_16_io_out_stage)
  );
  PE_1 local_pes_5_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_17_clock),
    .reset(local_pes_5_17_reset),
    .io_in_q(local_pes_5_17_io_in_q),
    .io_in_sum(local_pes_5_17_io_in_sum),
    .io_in_sum_exp(local_pes_5_17_io_in_sum_exp),
    .io_in_kv(local_pes_5_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_17_io_in_inv_sum),
    .io_in_stage(local_pes_5_17_io_in_stage),
    .io_out_q(local_pes_5_17_io_out_q),
    .io_out_sum(local_pes_5_17_io_out_sum),
    .io_out_sum_exp(local_pes_5_17_io_out_sum_exp),
    .io_out_kv(local_pes_5_17_io_out_kv),
    .io_out_stage(local_pes_5_17_io_out_stage)
  );
  PE_1 local_pes_5_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_18_clock),
    .reset(local_pes_5_18_reset),
    .io_in_q(local_pes_5_18_io_in_q),
    .io_in_sum(local_pes_5_18_io_in_sum),
    .io_in_sum_exp(local_pes_5_18_io_in_sum_exp),
    .io_in_kv(local_pes_5_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_18_io_in_inv_sum),
    .io_in_stage(local_pes_5_18_io_in_stage),
    .io_out_q(local_pes_5_18_io_out_q),
    .io_out_sum(local_pes_5_18_io_out_sum),
    .io_out_sum_exp(local_pes_5_18_io_out_sum_exp),
    .io_out_kv(local_pes_5_18_io_out_kv),
    .io_out_stage(local_pes_5_18_io_out_stage)
  );
  PE_1 local_pes_5_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_19_clock),
    .reset(local_pes_5_19_reset),
    .io_in_q(local_pes_5_19_io_in_q),
    .io_in_sum(local_pes_5_19_io_in_sum),
    .io_in_sum_exp(local_pes_5_19_io_in_sum_exp),
    .io_in_kv(local_pes_5_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_19_io_in_inv_sum),
    .io_in_stage(local_pes_5_19_io_in_stage),
    .io_out_q(local_pes_5_19_io_out_q),
    .io_out_sum(local_pes_5_19_io_out_sum),
    .io_out_sum_exp(local_pes_5_19_io_out_sum_exp),
    .io_out_kv(local_pes_5_19_io_out_kv),
    .io_out_stage(local_pes_5_19_io_out_stage)
  );
  PE_1 local_pes_5_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_20_clock),
    .reset(local_pes_5_20_reset),
    .io_in_q(local_pes_5_20_io_in_q),
    .io_in_sum(local_pes_5_20_io_in_sum),
    .io_in_sum_exp(local_pes_5_20_io_in_sum_exp),
    .io_in_kv(local_pes_5_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_20_io_in_inv_sum),
    .io_in_stage(local_pes_5_20_io_in_stage),
    .io_out_q(local_pes_5_20_io_out_q),
    .io_out_sum(local_pes_5_20_io_out_sum),
    .io_out_sum_exp(local_pes_5_20_io_out_sum_exp),
    .io_out_kv(local_pes_5_20_io_out_kv),
    .io_out_stage(local_pes_5_20_io_out_stage)
  );
  PE_1 local_pes_5_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_21_clock),
    .reset(local_pes_5_21_reset),
    .io_in_q(local_pes_5_21_io_in_q),
    .io_in_sum(local_pes_5_21_io_in_sum),
    .io_in_sum_exp(local_pes_5_21_io_in_sum_exp),
    .io_in_kv(local_pes_5_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_21_io_in_inv_sum),
    .io_in_stage(local_pes_5_21_io_in_stage),
    .io_out_q(local_pes_5_21_io_out_q),
    .io_out_sum(local_pes_5_21_io_out_sum),
    .io_out_sum_exp(local_pes_5_21_io_out_sum_exp),
    .io_out_kv(local_pes_5_21_io_out_kv),
    .io_out_stage(local_pes_5_21_io_out_stage)
  );
  PE_1 local_pes_5_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_22_clock),
    .reset(local_pes_5_22_reset),
    .io_in_q(local_pes_5_22_io_in_q),
    .io_in_sum(local_pes_5_22_io_in_sum),
    .io_in_sum_exp(local_pes_5_22_io_in_sum_exp),
    .io_in_kv(local_pes_5_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_22_io_in_inv_sum),
    .io_in_stage(local_pes_5_22_io_in_stage),
    .io_out_q(local_pes_5_22_io_out_q),
    .io_out_sum(local_pes_5_22_io_out_sum),
    .io_out_sum_exp(local_pes_5_22_io_out_sum_exp),
    .io_out_kv(local_pes_5_22_io_out_kv),
    .io_out_stage(local_pes_5_22_io_out_stage)
  );
  PE_1 local_pes_5_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_23_clock),
    .reset(local_pes_5_23_reset),
    .io_in_q(local_pes_5_23_io_in_q),
    .io_in_sum(local_pes_5_23_io_in_sum),
    .io_in_sum_exp(local_pes_5_23_io_in_sum_exp),
    .io_in_kv(local_pes_5_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_23_io_in_inv_sum),
    .io_in_stage(local_pes_5_23_io_in_stage),
    .io_out_q(local_pes_5_23_io_out_q),
    .io_out_sum(local_pes_5_23_io_out_sum),
    .io_out_sum_exp(local_pes_5_23_io_out_sum_exp),
    .io_out_kv(local_pes_5_23_io_out_kv),
    .io_out_stage(local_pes_5_23_io_out_stage)
  );
  PE_1 local_pes_5_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_24_clock),
    .reset(local_pes_5_24_reset),
    .io_in_q(local_pes_5_24_io_in_q),
    .io_in_sum(local_pes_5_24_io_in_sum),
    .io_in_sum_exp(local_pes_5_24_io_in_sum_exp),
    .io_in_kv(local_pes_5_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_24_io_in_inv_sum),
    .io_in_stage(local_pes_5_24_io_in_stage),
    .io_out_q(local_pes_5_24_io_out_q),
    .io_out_sum(local_pes_5_24_io_out_sum),
    .io_out_sum_exp(local_pes_5_24_io_out_sum_exp),
    .io_out_kv(local_pes_5_24_io_out_kv),
    .io_out_stage(local_pes_5_24_io_out_stage)
  );
  PE_1 local_pes_5_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_25_clock),
    .reset(local_pes_5_25_reset),
    .io_in_q(local_pes_5_25_io_in_q),
    .io_in_sum(local_pes_5_25_io_in_sum),
    .io_in_sum_exp(local_pes_5_25_io_in_sum_exp),
    .io_in_kv(local_pes_5_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_25_io_in_inv_sum),
    .io_in_stage(local_pes_5_25_io_in_stage),
    .io_out_q(local_pes_5_25_io_out_q),
    .io_out_sum(local_pes_5_25_io_out_sum),
    .io_out_sum_exp(local_pes_5_25_io_out_sum_exp),
    .io_out_kv(local_pes_5_25_io_out_kv),
    .io_out_stage(local_pes_5_25_io_out_stage)
  );
  PE_1 local_pes_5_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_26_clock),
    .reset(local_pes_5_26_reset),
    .io_in_q(local_pes_5_26_io_in_q),
    .io_in_sum(local_pes_5_26_io_in_sum),
    .io_in_sum_exp(local_pes_5_26_io_in_sum_exp),
    .io_in_kv(local_pes_5_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_26_io_in_inv_sum),
    .io_in_stage(local_pes_5_26_io_in_stage),
    .io_out_q(local_pes_5_26_io_out_q),
    .io_out_sum(local_pes_5_26_io_out_sum),
    .io_out_sum_exp(local_pes_5_26_io_out_sum_exp),
    .io_out_kv(local_pes_5_26_io_out_kv),
    .io_out_stage(local_pes_5_26_io_out_stage)
  );
  PE_1 local_pes_5_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_27_clock),
    .reset(local_pes_5_27_reset),
    .io_in_q(local_pes_5_27_io_in_q),
    .io_in_sum(local_pes_5_27_io_in_sum),
    .io_in_sum_exp(local_pes_5_27_io_in_sum_exp),
    .io_in_kv(local_pes_5_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_27_io_in_inv_sum),
    .io_in_stage(local_pes_5_27_io_in_stage),
    .io_out_q(local_pes_5_27_io_out_q),
    .io_out_sum(local_pes_5_27_io_out_sum),
    .io_out_sum_exp(local_pes_5_27_io_out_sum_exp),
    .io_out_kv(local_pes_5_27_io_out_kv),
    .io_out_stage(local_pes_5_27_io_out_stage)
  );
  PE_1 local_pes_5_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_28_clock),
    .reset(local_pes_5_28_reset),
    .io_in_q(local_pes_5_28_io_in_q),
    .io_in_sum(local_pes_5_28_io_in_sum),
    .io_in_sum_exp(local_pes_5_28_io_in_sum_exp),
    .io_in_kv(local_pes_5_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_28_io_in_inv_sum),
    .io_in_stage(local_pes_5_28_io_in_stage),
    .io_out_q(local_pes_5_28_io_out_q),
    .io_out_sum(local_pes_5_28_io_out_sum),
    .io_out_sum_exp(local_pes_5_28_io_out_sum_exp),
    .io_out_kv(local_pes_5_28_io_out_kv),
    .io_out_stage(local_pes_5_28_io_out_stage)
  );
  PE_1 local_pes_5_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_29_clock),
    .reset(local_pes_5_29_reset),
    .io_in_q(local_pes_5_29_io_in_q),
    .io_in_sum(local_pes_5_29_io_in_sum),
    .io_in_sum_exp(local_pes_5_29_io_in_sum_exp),
    .io_in_kv(local_pes_5_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_29_io_in_inv_sum),
    .io_in_stage(local_pes_5_29_io_in_stage),
    .io_out_q(local_pes_5_29_io_out_q),
    .io_out_sum(local_pes_5_29_io_out_sum),
    .io_out_sum_exp(local_pes_5_29_io_out_sum_exp),
    .io_out_kv(local_pes_5_29_io_out_kv),
    .io_out_stage(local_pes_5_29_io_out_stage)
  );
  PE_1 local_pes_5_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_30_clock),
    .reset(local_pes_5_30_reset),
    .io_in_q(local_pes_5_30_io_in_q),
    .io_in_sum(local_pes_5_30_io_in_sum),
    .io_in_sum_exp(local_pes_5_30_io_in_sum_exp),
    .io_in_kv(local_pes_5_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_30_io_in_inv_sum),
    .io_in_stage(local_pes_5_30_io_in_stage),
    .io_out_q(local_pes_5_30_io_out_q),
    .io_out_sum(local_pes_5_30_io_out_sum),
    .io_out_sum_exp(local_pes_5_30_io_out_sum_exp),
    .io_out_kv(local_pes_5_30_io_out_kv),
    .io_out_stage(local_pes_5_30_io_out_stage)
  );
  PE_1 local_pes_5_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_5_31_clock),
    .reset(local_pes_5_31_reset),
    .io_in_q(local_pes_5_31_io_in_q),
    .io_in_sum(local_pes_5_31_io_in_sum),
    .io_in_sum_exp(local_pes_5_31_io_in_sum_exp),
    .io_in_kv(local_pes_5_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_5_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_5_31_io_in_inv_sum),
    .io_in_stage(local_pes_5_31_io_in_stage),
    .io_out_q(local_pes_5_31_io_out_q),
    .io_out_sum(local_pes_5_31_io_out_sum),
    .io_out_sum_exp(local_pes_5_31_io_out_sum_exp),
    .io_out_kv(local_pes_5_31_io_out_kv),
    .io_out_stage(local_pes_5_31_io_out_stage)
  );
  PE local_pes_6_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_0_clock),
    .reset(local_pes_6_0_reset),
    .io_in_q(local_pes_6_0_io_in_q),
    .io_in_kv(local_pes_6_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_0_io_in_inv_sum),
    .io_in_stage(local_pes_6_0_io_in_stage),
    .io_out_q(local_pes_6_0_io_out_q),
    .io_out_sum(local_pes_6_0_io_out_sum),
    .io_out_kv(local_pes_6_0_io_out_kv),
    .io_out_stage(local_pes_6_0_io_out_stage)
  );
  PE_1 local_pes_6_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_1_clock),
    .reset(local_pes_6_1_reset),
    .io_in_q(local_pes_6_1_io_in_q),
    .io_in_sum(local_pes_6_1_io_in_sum),
    .io_in_sum_exp(local_pes_6_1_io_in_sum_exp),
    .io_in_kv(local_pes_6_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_1_io_in_inv_sum),
    .io_in_stage(local_pes_6_1_io_in_stage),
    .io_out_q(local_pes_6_1_io_out_q),
    .io_out_sum(local_pes_6_1_io_out_sum),
    .io_out_sum_exp(local_pes_6_1_io_out_sum_exp),
    .io_out_kv(local_pes_6_1_io_out_kv),
    .io_out_stage(local_pes_6_1_io_out_stage)
  );
  PE_1 local_pes_6_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_2_clock),
    .reset(local_pes_6_2_reset),
    .io_in_q(local_pes_6_2_io_in_q),
    .io_in_sum(local_pes_6_2_io_in_sum),
    .io_in_sum_exp(local_pes_6_2_io_in_sum_exp),
    .io_in_kv(local_pes_6_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_2_io_in_inv_sum),
    .io_in_stage(local_pes_6_2_io_in_stage),
    .io_out_q(local_pes_6_2_io_out_q),
    .io_out_sum(local_pes_6_2_io_out_sum),
    .io_out_sum_exp(local_pes_6_2_io_out_sum_exp),
    .io_out_kv(local_pes_6_2_io_out_kv),
    .io_out_stage(local_pes_6_2_io_out_stage)
  );
  PE_1 local_pes_6_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_3_clock),
    .reset(local_pes_6_3_reset),
    .io_in_q(local_pes_6_3_io_in_q),
    .io_in_sum(local_pes_6_3_io_in_sum),
    .io_in_sum_exp(local_pes_6_3_io_in_sum_exp),
    .io_in_kv(local_pes_6_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_3_io_in_inv_sum),
    .io_in_stage(local_pes_6_3_io_in_stage),
    .io_out_q(local_pes_6_3_io_out_q),
    .io_out_sum(local_pes_6_3_io_out_sum),
    .io_out_sum_exp(local_pes_6_3_io_out_sum_exp),
    .io_out_kv(local_pes_6_3_io_out_kv),
    .io_out_stage(local_pes_6_3_io_out_stage)
  );
  PE_1 local_pes_6_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_4_clock),
    .reset(local_pes_6_4_reset),
    .io_in_q(local_pes_6_4_io_in_q),
    .io_in_sum(local_pes_6_4_io_in_sum),
    .io_in_sum_exp(local_pes_6_4_io_in_sum_exp),
    .io_in_kv(local_pes_6_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_4_io_in_inv_sum),
    .io_in_stage(local_pes_6_4_io_in_stage),
    .io_out_q(local_pes_6_4_io_out_q),
    .io_out_sum(local_pes_6_4_io_out_sum),
    .io_out_sum_exp(local_pes_6_4_io_out_sum_exp),
    .io_out_kv(local_pes_6_4_io_out_kv),
    .io_out_stage(local_pes_6_4_io_out_stage)
  );
  PE_1 local_pes_6_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_5_clock),
    .reset(local_pes_6_5_reset),
    .io_in_q(local_pes_6_5_io_in_q),
    .io_in_sum(local_pes_6_5_io_in_sum),
    .io_in_sum_exp(local_pes_6_5_io_in_sum_exp),
    .io_in_kv(local_pes_6_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_5_io_in_inv_sum),
    .io_in_stage(local_pes_6_5_io_in_stage),
    .io_out_q(local_pes_6_5_io_out_q),
    .io_out_sum(local_pes_6_5_io_out_sum),
    .io_out_sum_exp(local_pes_6_5_io_out_sum_exp),
    .io_out_kv(local_pes_6_5_io_out_kv),
    .io_out_stage(local_pes_6_5_io_out_stage)
  );
  PE_1 local_pes_6_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_6_clock),
    .reset(local_pes_6_6_reset),
    .io_in_q(local_pes_6_6_io_in_q),
    .io_in_sum(local_pes_6_6_io_in_sum),
    .io_in_sum_exp(local_pes_6_6_io_in_sum_exp),
    .io_in_kv(local_pes_6_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_6_io_in_inv_sum),
    .io_in_stage(local_pes_6_6_io_in_stage),
    .io_out_q(local_pes_6_6_io_out_q),
    .io_out_sum(local_pes_6_6_io_out_sum),
    .io_out_sum_exp(local_pes_6_6_io_out_sum_exp),
    .io_out_kv(local_pes_6_6_io_out_kv),
    .io_out_stage(local_pes_6_6_io_out_stage)
  );
  PE_1 local_pes_6_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_7_clock),
    .reset(local_pes_6_7_reset),
    .io_in_q(local_pes_6_7_io_in_q),
    .io_in_sum(local_pes_6_7_io_in_sum),
    .io_in_sum_exp(local_pes_6_7_io_in_sum_exp),
    .io_in_kv(local_pes_6_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_7_io_in_inv_sum),
    .io_in_stage(local_pes_6_7_io_in_stage),
    .io_out_q(local_pes_6_7_io_out_q),
    .io_out_sum(local_pes_6_7_io_out_sum),
    .io_out_sum_exp(local_pes_6_7_io_out_sum_exp),
    .io_out_kv(local_pes_6_7_io_out_kv),
    .io_out_stage(local_pes_6_7_io_out_stage)
  );
  PE_1 local_pes_6_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_8_clock),
    .reset(local_pes_6_8_reset),
    .io_in_q(local_pes_6_8_io_in_q),
    .io_in_sum(local_pes_6_8_io_in_sum),
    .io_in_sum_exp(local_pes_6_8_io_in_sum_exp),
    .io_in_kv(local_pes_6_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_8_io_in_inv_sum),
    .io_in_stage(local_pes_6_8_io_in_stage),
    .io_out_q(local_pes_6_8_io_out_q),
    .io_out_sum(local_pes_6_8_io_out_sum),
    .io_out_sum_exp(local_pes_6_8_io_out_sum_exp),
    .io_out_kv(local_pes_6_8_io_out_kv),
    .io_out_stage(local_pes_6_8_io_out_stage)
  );
  PE_1 local_pes_6_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_9_clock),
    .reset(local_pes_6_9_reset),
    .io_in_q(local_pes_6_9_io_in_q),
    .io_in_sum(local_pes_6_9_io_in_sum),
    .io_in_sum_exp(local_pes_6_9_io_in_sum_exp),
    .io_in_kv(local_pes_6_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_9_io_in_inv_sum),
    .io_in_stage(local_pes_6_9_io_in_stage),
    .io_out_q(local_pes_6_9_io_out_q),
    .io_out_sum(local_pes_6_9_io_out_sum),
    .io_out_sum_exp(local_pes_6_9_io_out_sum_exp),
    .io_out_kv(local_pes_6_9_io_out_kv),
    .io_out_stage(local_pes_6_9_io_out_stage)
  );
  PE_1 local_pes_6_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_10_clock),
    .reset(local_pes_6_10_reset),
    .io_in_q(local_pes_6_10_io_in_q),
    .io_in_sum(local_pes_6_10_io_in_sum),
    .io_in_sum_exp(local_pes_6_10_io_in_sum_exp),
    .io_in_kv(local_pes_6_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_10_io_in_inv_sum),
    .io_in_stage(local_pes_6_10_io_in_stage),
    .io_out_q(local_pes_6_10_io_out_q),
    .io_out_sum(local_pes_6_10_io_out_sum),
    .io_out_sum_exp(local_pes_6_10_io_out_sum_exp),
    .io_out_kv(local_pes_6_10_io_out_kv),
    .io_out_stage(local_pes_6_10_io_out_stage)
  );
  PE_1 local_pes_6_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_11_clock),
    .reset(local_pes_6_11_reset),
    .io_in_q(local_pes_6_11_io_in_q),
    .io_in_sum(local_pes_6_11_io_in_sum),
    .io_in_sum_exp(local_pes_6_11_io_in_sum_exp),
    .io_in_kv(local_pes_6_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_11_io_in_inv_sum),
    .io_in_stage(local_pes_6_11_io_in_stage),
    .io_out_q(local_pes_6_11_io_out_q),
    .io_out_sum(local_pes_6_11_io_out_sum),
    .io_out_sum_exp(local_pes_6_11_io_out_sum_exp),
    .io_out_kv(local_pes_6_11_io_out_kv),
    .io_out_stage(local_pes_6_11_io_out_stage)
  );
  PE_1 local_pes_6_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_12_clock),
    .reset(local_pes_6_12_reset),
    .io_in_q(local_pes_6_12_io_in_q),
    .io_in_sum(local_pes_6_12_io_in_sum),
    .io_in_sum_exp(local_pes_6_12_io_in_sum_exp),
    .io_in_kv(local_pes_6_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_12_io_in_inv_sum),
    .io_in_stage(local_pes_6_12_io_in_stage),
    .io_out_q(local_pes_6_12_io_out_q),
    .io_out_sum(local_pes_6_12_io_out_sum),
    .io_out_sum_exp(local_pes_6_12_io_out_sum_exp),
    .io_out_kv(local_pes_6_12_io_out_kv),
    .io_out_stage(local_pes_6_12_io_out_stage)
  );
  PE_1 local_pes_6_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_13_clock),
    .reset(local_pes_6_13_reset),
    .io_in_q(local_pes_6_13_io_in_q),
    .io_in_sum(local_pes_6_13_io_in_sum),
    .io_in_sum_exp(local_pes_6_13_io_in_sum_exp),
    .io_in_kv(local_pes_6_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_13_io_in_inv_sum),
    .io_in_stage(local_pes_6_13_io_in_stage),
    .io_out_q(local_pes_6_13_io_out_q),
    .io_out_sum(local_pes_6_13_io_out_sum),
    .io_out_sum_exp(local_pes_6_13_io_out_sum_exp),
    .io_out_kv(local_pes_6_13_io_out_kv),
    .io_out_stage(local_pes_6_13_io_out_stage)
  );
  PE_1 local_pes_6_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_14_clock),
    .reset(local_pes_6_14_reset),
    .io_in_q(local_pes_6_14_io_in_q),
    .io_in_sum(local_pes_6_14_io_in_sum),
    .io_in_sum_exp(local_pes_6_14_io_in_sum_exp),
    .io_in_kv(local_pes_6_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_14_io_in_inv_sum),
    .io_in_stage(local_pes_6_14_io_in_stage),
    .io_out_q(local_pes_6_14_io_out_q),
    .io_out_sum(local_pes_6_14_io_out_sum),
    .io_out_sum_exp(local_pes_6_14_io_out_sum_exp),
    .io_out_kv(local_pes_6_14_io_out_kv),
    .io_out_stage(local_pes_6_14_io_out_stage)
  );
  PE_1 local_pes_6_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_15_clock),
    .reset(local_pes_6_15_reset),
    .io_in_q(local_pes_6_15_io_in_q),
    .io_in_sum(local_pes_6_15_io_in_sum),
    .io_in_sum_exp(local_pes_6_15_io_in_sum_exp),
    .io_in_kv(local_pes_6_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_15_io_in_inv_sum),
    .io_in_stage(local_pes_6_15_io_in_stage),
    .io_out_q(local_pes_6_15_io_out_q),
    .io_out_sum(local_pes_6_15_io_out_sum),
    .io_out_sum_exp(local_pes_6_15_io_out_sum_exp),
    .io_out_kv(local_pes_6_15_io_out_kv),
    .io_out_stage(local_pes_6_15_io_out_stage)
  );
  PE_1 local_pes_6_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_16_clock),
    .reset(local_pes_6_16_reset),
    .io_in_q(local_pes_6_16_io_in_q),
    .io_in_sum(local_pes_6_16_io_in_sum),
    .io_in_sum_exp(local_pes_6_16_io_in_sum_exp),
    .io_in_kv(local_pes_6_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_16_io_in_inv_sum),
    .io_in_stage(local_pes_6_16_io_in_stage),
    .io_out_q(local_pes_6_16_io_out_q),
    .io_out_sum(local_pes_6_16_io_out_sum),
    .io_out_sum_exp(local_pes_6_16_io_out_sum_exp),
    .io_out_kv(local_pes_6_16_io_out_kv),
    .io_out_stage(local_pes_6_16_io_out_stage)
  );
  PE_1 local_pes_6_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_17_clock),
    .reset(local_pes_6_17_reset),
    .io_in_q(local_pes_6_17_io_in_q),
    .io_in_sum(local_pes_6_17_io_in_sum),
    .io_in_sum_exp(local_pes_6_17_io_in_sum_exp),
    .io_in_kv(local_pes_6_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_17_io_in_inv_sum),
    .io_in_stage(local_pes_6_17_io_in_stage),
    .io_out_q(local_pes_6_17_io_out_q),
    .io_out_sum(local_pes_6_17_io_out_sum),
    .io_out_sum_exp(local_pes_6_17_io_out_sum_exp),
    .io_out_kv(local_pes_6_17_io_out_kv),
    .io_out_stage(local_pes_6_17_io_out_stage)
  );
  PE_1 local_pes_6_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_18_clock),
    .reset(local_pes_6_18_reset),
    .io_in_q(local_pes_6_18_io_in_q),
    .io_in_sum(local_pes_6_18_io_in_sum),
    .io_in_sum_exp(local_pes_6_18_io_in_sum_exp),
    .io_in_kv(local_pes_6_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_18_io_in_inv_sum),
    .io_in_stage(local_pes_6_18_io_in_stage),
    .io_out_q(local_pes_6_18_io_out_q),
    .io_out_sum(local_pes_6_18_io_out_sum),
    .io_out_sum_exp(local_pes_6_18_io_out_sum_exp),
    .io_out_kv(local_pes_6_18_io_out_kv),
    .io_out_stage(local_pes_6_18_io_out_stage)
  );
  PE_1 local_pes_6_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_19_clock),
    .reset(local_pes_6_19_reset),
    .io_in_q(local_pes_6_19_io_in_q),
    .io_in_sum(local_pes_6_19_io_in_sum),
    .io_in_sum_exp(local_pes_6_19_io_in_sum_exp),
    .io_in_kv(local_pes_6_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_19_io_in_inv_sum),
    .io_in_stage(local_pes_6_19_io_in_stage),
    .io_out_q(local_pes_6_19_io_out_q),
    .io_out_sum(local_pes_6_19_io_out_sum),
    .io_out_sum_exp(local_pes_6_19_io_out_sum_exp),
    .io_out_kv(local_pes_6_19_io_out_kv),
    .io_out_stage(local_pes_6_19_io_out_stage)
  );
  PE_1 local_pes_6_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_20_clock),
    .reset(local_pes_6_20_reset),
    .io_in_q(local_pes_6_20_io_in_q),
    .io_in_sum(local_pes_6_20_io_in_sum),
    .io_in_sum_exp(local_pes_6_20_io_in_sum_exp),
    .io_in_kv(local_pes_6_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_20_io_in_inv_sum),
    .io_in_stage(local_pes_6_20_io_in_stage),
    .io_out_q(local_pes_6_20_io_out_q),
    .io_out_sum(local_pes_6_20_io_out_sum),
    .io_out_sum_exp(local_pes_6_20_io_out_sum_exp),
    .io_out_kv(local_pes_6_20_io_out_kv),
    .io_out_stage(local_pes_6_20_io_out_stage)
  );
  PE_1 local_pes_6_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_21_clock),
    .reset(local_pes_6_21_reset),
    .io_in_q(local_pes_6_21_io_in_q),
    .io_in_sum(local_pes_6_21_io_in_sum),
    .io_in_sum_exp(local_pes_6_21_io_in_sum_exp),
    .io_in_kv(local_pes_6_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_21_io_in_inv_sum),
    .io_in_stage(local_pes_6_21_io_in_stage),
    .io_out_q(local_pes_6_21_io_out_q),
    .io_out_sum(local_pes_6_21_io_out_sum),
    .io_out_sum_exp(local_pes_6_21_io_out_sum_exp),
    .io_out_kv(local_pes_6_21_io_out_kv),
    .io_out_stage(local_pes_6_21_io_out_stage)
  );
  PE_1 local_pes_6_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_22_clock),
    .reset(local_pes_6_22_reset),
    .io_in_q(local_pes_6_22_io_in_q),
    .io_in_sum(local_pes_6_22_io_in_sum),
    .io_in_sum_exp(local_pes_6_22_io_in_sum_exp),
    .io_in_kv(local_pes_6_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_22_io_in_inv_sum),
    .io_in_stage(local_pes_6_22_io_in_stage),
    .io_out_q(local_pes_6_22_io_out_q),
    .io_out_sum(local_pes_6_22_io_out_sum),
    .io_out_sum_exp(local_pes_6_22_io_out_sum_exp),
    .io_out_kv(local_pes_6_22_io_out_kv),
    .io_out_stage(local_pes_6_22_io_out_stage)
  );
  PE_1 local_pes_6_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_23_clock),
    .reset(local_pes_6_23_reset),
    .io_in_q(local_pes_6_23_io_in_q),
    .io_in_sum(local_pes_6_23_io_in_sum),
    .io_in_sum_exp(local_pes_6_23_io_in_sum_exp),
    .io_in_kv(local_pes_6_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_23_io_in_inv_sum),
    .io_in_stage(local_pes_6_23_io_in_stage),
    .io_out_q(local_pes_6_23_io_out_q),
    .io_out_sum(local_pes_6_23_io_out_sum),
    .io_out_sum_exp(local_pes_6_23_io_out_sum_exp),
    .io_out_kv(local_pes_6_23_io_out_kv),
    .io_out_stage(local_pes_6_23_io_out_stage)
  );
  PE_1 local_pes_6_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_24_clock),
    .reset(local_pes_6_24_reset),
    .io_in_q(local_pes_6_24_io_in_q),
    .io_in_sum(local_pes_6_24_io_in_sum),
    .io_in_sum_exp(local_pes_6_24_io_in_sum_exp),
    .io_in_kv(local_pes_6_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_24_io_in_inv_sum),
    .io_in_stage(local_pes_6_24_io_in_stage),
    .io_out_q(local_pes_6_24_io_out_q),
    .io_out_sum(local_pes_6_24_io_out_sum),
    .io_out_sum_exp(local_pes_6_24_io_out_sum_exp),
    .io_out_kv(local_pes_6_24_io_out_kv),
    .io_out_stage(local_pes_6_24_io_out_stage)
  );
  PE_1 local_pes_6_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_25_clock),
    .reset(local_pes_6_25_reset),
    .io_in_q(local_pes_6_25_io_in_q),
    .io_in_sum(local_pes_6_25_io_in_sum),
    .io_in_sum_exp(local_pes_6_25_io_in_sum_exp),
    .io_in_kv(local_pes_6_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_25_io_in_inv_sum),
    .io_in_stage(local_pes_6_25_io_in_stage),
    .io_out_q(local_pes_6_25_io_out_q),
    .io_out_sum(local_pes_6_25_io_out_sum),
    .io_out_sum_exp(local_pes_6_25_io_out_sum_exp),
    .io_out_kv(local_pes_6_25_io_out_kv),
    .io_out_stage(local_pes_6_25_io_out_stage)
  );
  PE_1 local_pes_6_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_26_clock),
    .reset(local_pes_6_26_reset),
    .io_in_q(local_pes_6_26_io_in_q),
    .io_in_sum(local_pes_6_26_io_in_sum),
    .io_in_sum_exp(local_pes_6_26_io_in_sum_exp),
    .io_in_kv(local_pes_6_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_26_io_in_inv_sum),
    .io_in_stage(local_pes_6_26_io_in_stage),
    .io_out_q(local_pes_6_26_io_out_q),
    .io_out_sum(local_pes_6_26_io_out_sum),
    .io_out_sum_exp(local_pes_6_26_io_out_sum_exp),
    .io_out_kv(local_pes_6_26_io_out_kv),
    .io_out_stage(local_pes_6_26_io_out_stage)
  );
  PE_1 local_pes_6_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_27_clock),
    .reset(local_pes_6_27_reset),
    .io_in_q(local_pes_6_27_io_in_q),
    .io_in_sum(local_pes_6_27_io_in_sum),
    .io_in_sum_exp(local_pes_6_27_io_in_sum_exp),
    .io_in_kv(local_pes_6_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_27_io_in_inv_sum),
    .io_in_stage(local_pes_6_27_io_in_stage),
    .io_out_q(local_pes_6_27_io_out_q),
    .io_out_sum(local_pes_6_27_io_out_sum),
    .io_out_sum_exp(local_pes_6_27_io_out_sum_exp),
    .io_out_kv(local_pes_6_27_io_out_kv),
    .io_out_stage(local_pes_6_27_io_out_stage)
  );
  PE_1 local_pes_6_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_28_clock),
    .reset(local_pes_6_28_reset),
    .io_in_q(local_pes_6_28_io_in_q),
    .io_in_sum(local_pes_6_28_io_in_sum),
    .io_in_sum_exp(local_pes_6_28_io_in_sum_exp),
    .io_in_kv(local_pes_6_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_28_io_in_inv_sum),
    .io_in_stage(local_pes_6_28_io_in_stage),
    .io_out_q(local_pes_6_28_io_out_q),
    .io_out_sum(local_pes_6_28_io_out_sum),
    .io_out_sum_exp(local_pes_6_28_io_out_sum_exp),
    .io_out_kv(local_pes_6_28_io_out_kv),
    .io_out_stage(local_pes_6_28_io_out_stage)
  );
  PE_1 local_pes_6_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_29_clock),
    .reset(local_pes_6_29_reset),
    .io_in_q(local_pes_6_29_io_in_q),
    .io_in_sum(local_pes_6_29_io_in_sum),
    .io_in_sum_exp(local_pes_6_29_io_in_sum_exp),
    .io_in_kv(local_pes_6_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_29_io_in_inv_sum),
    .io_in_stage(local_pes_6_29_io_in_stage),
    .io_out_q(local_pes_6_29_io_out_q),
    .io_out_sum(local_pes_6_29_io_out_sum),
    .io_out_sum_exp(local_pes_6_29_io_out_sum_exp),
    .io_out_kv(local_pes_6_29_io_out_kv),
    .io_out_stage(local_pes_6_29_io_out_stage)
  );
  PE_1 local_pes_6_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_30_clock),
    .reset(local_pes_6_30_reset),
    .io_in_q(local_pes_6_30_io_in_q),
    .io_in_sum(local_pes_6_30_io_in_sum),
    .io_in_sum_exp(local_pes_6_30_io_in_sum_exp),
    .io_in_kv(local_pes_6_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_30_io_in_inv_sum),
    .io_in_stage(local_pes_6_30_io_in_stage),
    .io_out_q(local_pes_6_30_io_out_q),
    .io_out_sum(local_pes_6_30_io_out_sum),
    .io_out_sum_exp(local_pes_6_30_io_out_sum_exp),
    .io_out_kv(local_pes_6_30_io_out_kv),
    .io_out_stage(local_pes_6_30_io_out_stage)
  );
  PE_1 local_pes_6_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_6_31_clock),
    .reset(local_pes_6_31_reset),
    .io_in_q(local_pes_6_31_io_in_q),
    .io_in_sum(local_pes_6_31_io_in_sum),
    .io_in_sum_exp(local_pes_6_31_io_in_sum_exp),
    .io_in_kv(local_pes_6_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_6_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_6_31_io_in_inv_sum),
    .io_in_stage(local_pes_6_31_io_in_stage),
    .io_out_q(local_pes_6_31_io_out_q),
    .io_out_sum(local_pes_6_31_io_out_sum),
    .io_out_sum_exp(local_pes_6_31_io_out_sum_exp),
    .io_out_kv(local_pes_6_31_io_out_kv),
    .io_out_stage(local_pes_6_31_io_out_stage)
  );
  PE local_pes_7_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_0_clock),
    .reset(local_pes_7_0_reset),
    .io_in_q(local_pes_7_0_io_in_q),
    .io_in_kv(local_pes_7_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_0_io_in_inv_sum),
    .io_in_stage(local_pes_7_0_io_in_stage),
    .io_out_q(local_pes_7_0_io_out_q),
    .io_out_sum(local_pes_7_0_io_out_sum),
    .io_out_kv(local_pes_7_0_io_out_kv),
    .io_out_stage(local_pes_7_0_io_out_stage)
  );
  PE_1 local_pes_7_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_1_clock),
    .reset(local_pes_7_1_reset),
    .io_in_q(local_pes_7_1_io_in_q),
    .io_in_sum(local_pes_7_1_io_in_sum),
    .io_in_sum_exp(local_pes_7_1_io_in_sum_exp),
    .io_in_kv(local_pes_7_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_1_io_in_inv_sum),
    .io_in_stage(local_pes_7_1_io_in_stage),
    .io_out_q(local_pes_7_1_io_out_q),
    .io_out_sum(local_pes_7_1_io_out_sum),
    .io_out_sum_exp(local_pes_7_1_io_out_sum_exp),
    .io_out_kv(local_pes_7_1_io_out_kv),
    .io_out_stage(local_pes_7_1_io_out_stage)
  );
  PE_1 local_pes_7_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_2_clock),
    .reset(local_pes_7_2_reset),
    .io_in_q(local_pes_7_2_io_in_q),
    .io_in_sum(local_pes_7_2_io_in_sum),
    .io_in_sum_exp(local_pes_7_2_io_in_sum_exp),
    .io_in_kv(local_pes_7_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_2_io_in_inv_sum),
    .io_in_stage(local_pes_7_2_io_in_stage),
    .io_out_q(local_pes_7_2_io_out_q),
    .io_out_sum(local_pes_7_2_io_out_sum),
    .io_out_sum_exp(local_pes_7_2_io_out_sum_exp),
    .io_out_kv(local_pes_7_2_io_out_kv),
    .io_out_stage(local_pes_7_2_io_out_stage)
  );
  PE_1 local_pes_7_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_3_clock),
    .reset(local_pes_7_3_reset),
    .io_in_q(local_pes_7_3_io_in_q),
    .io_in_sum(local_pes_7_3_io_in_sum),
    .io_in_sum_exp(local_pes_7_3_io_in_sum_exp),
    .io_in_kv(local_pes_7_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_3_io_in_inv_sum),
    .io_in_stage(local_pes_7_3_io_in_stage),
    .io_out_q(local_pes_7_3_io_out_q),
    .io_out_sum(local_pes_7_3_io_out_sum),
    .io_out_sum_exp(local_pes_7_3_io_out_sum_exp),
    .io_out_kv(local_pes_7_3_io_out_kv),
    .io_out_stage(local_pes_7_3_io_out_stage)
  );
  PE_1 local_pes_7_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_4_clock),
    .reset(local_pes_7_4_reset),
    .io_in_q(local_pes_7_4_io_in_q),
    .io_in_sum(local_pes_7_4_io_in_sum),
    .io_in_sum_exp(local_pes_7_4_io_in_sum_exp),
    .io_in_kv(local_pes_7_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_4_io_in_inv_sum),
    .io_in_stage(local_pes_7_4_io_in_stage),
    .io_out_q(local_pes_7_4_io_out_q),
    .io_out_sum(local_pes_7_4_io_out_sum),
    .io_out_sum_exp(local_pes_7_4_io_out_sum_exp),
    .io_out_kv(local_pes_7_4_io_out_kv),
    .io_out_stage(local_pes_7_4_io_out_stage)
  );
  PE_1 local_pes_7_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_5_clock),
    .reset(local_pes_7_5_reset),
    .io_in_q(local_pes_7_5_io_in_q),
    .io_in_sum(local_pes_7_5_io_in_sum),
    .io_in_sum_exp(local_pes_7_5_io_in_sum_exp),
    .io_in_kv(local_pes_7_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_5_io_in_inv_sum),
    .io_in_stage(local_pes_7_5_io_in_stage),
    .io_out_q(local_pes_7_5_io_out_q),
    .io_out_sum(local_pes_7_5_io_out_sum),
    .io_out_sum_exp(local_pes_7_5_io_out_sum_exp),
    .io_out_kv(local_pes_7_5_io_out_kv),
    .io_out_stage(local_pes_7_5_io_out_stage)
  );
  PE_1 local_pes_7_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_6_clock),
    .reset(local_pes_7_6_reset),
    .io_in_q(local_pes_7_6_io_in_q),
    .io_in_sum(local_pes_7_6_io_in_sum),
    .io_in_sum_exp(local_pes_7_6_io_in_sum_exp),
    .io_in_kv(local_pes_7_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_6_io_in_inv_sum),
    .io_in_stage(local_pes_7_6_io_in_stage),
    .io_out_q(local_pes_7_6_io_out_q),
    .io_out_sum(local_pes_7_6_io_out_sum),
    .io_out_sum_exp(local_pes_7_6_io_out_sum_exp),
    .io_out_kv(local_pes_7_6_io_out_kv),
    .io_out_stage(local_pes_7_6_io_out_stage)
  );
  PE_1 local_pes_7_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_7_clock),
    .reset(local_pes_7_7_reset),
    .io_in_q(local_pes_7_7_io_in_q),
    .io_in_sum(local_pes_7_7_io_in_sum),
    .io_in_sum_exp(local_pes_7_7_io_in_sum_exp),
    .io_in_kv(local_pes_7_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_7_io_in_inv_sum),
    .io_in_stage(local_pes_7_7_io_in_stage),
    .io_out_q(local_pes_7_7_io_out_q),
    .io_out_sum(local_pes_7_7_io_out_sum),
    .io_out_sum_exp(local_pes_7_7_io_out_sum_exp),
    .io_out_kv(local_pes_7_7_io_out_kv),
    .io_out_stage(local_pes_7_7_io_out_stage)
  );
  PE_1 local_pes_7_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_8_clock),
    .reset(local_pes_7_8_reset),
    .io_in_q(local_pes_7_8_io_in_q),
    .io_in_sum(local_pes_7_8_io_in_sum),
    .io_in_sum_exp(local_pes_7_8_io_in_sum_exp),
    .io_in_kv(local_pes_7_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_8_io_in_inv_sum),
    .io_in_stage(local_pes_7_8_io_in_stage),
    .io_out_q(local_pes_7_8_io_out_q),
    .io_out_sum(local_pes_7_8_io_out_sum),
    .io_out_sum_exp(local_pes_7_8_io_out_sum_exp),
    .io_out_kv(local_pes_7_8_io_out_kv),
    .io_out_stage(local_pes_7_8_io_out_stage)
  );
  PE_1 local_pes_7_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_9_clock),
    .reset(local_pes_7_9_reset),
    .io_in_q(local_pes_7_9_io_in_q),
    .io_in_sum(local_pes_7_9_io_in_sum),
    .io_in_sum_exp(local_pes_7_9_io_in_sum_exp),
    .io_in_kv(local_pes_7_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_9_io_in_inv_sum),
    .io_in_stage(local_pes_7_9_io_in_stage),
    .io_out_q(local_pes_7_9_io_out_q),
    .io_out_sum(local_pes_7_9_io_out_sum),
    .io_out_sum_exp(local_pes_7_9_io_out_sum_exp),
    .io_out_kv(local_pes_7_9_io_out_kv),
    .io_out_stage(local_pes_7_9_io_out_stage)
  );
  PE_1 local_pes_7_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_10_clock),
    .reset(local_pes_7_10_reset),
    .io_in_q(local_pes_7_10_io_in_q),
    .io_in_sum(local_pes_7_10_io_in_sum),
    .io_in_sum_exp(local_pes_7_10_io_in_sum_exp),
    .io_in_kv(local_pes_7_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_10_io_in_inv_sum),
    .io_in_stage(local_pes_7_10_io_in_stage),
    .io_out_q(local_pes_7_10_io_out_q),
    .io_out_sum(local_pes_7_10_io_out_sum),
    .io_out_sum_exp(local_pes_7_10_io_out_sum_exp),
    .io_out_kv(local_pes_7_10_io_out_kv),
    .io_out_stage(local_pes_7_10_io_out_stage)
  );
  PE_1 local_pes_7_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_11_clock),
    .reset(local_pes_7_11_reset),
    .io_in_q(local_pes_7_11_io_in_q),
    .io_in_sum(local_pes_7_11_io_in_sum),
    .io_in_sum_exp(local_pes_7_11_io_in_sum_exp),
    .io_in_kv(local_pes_7_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_11_io_in_inv_sum),
    .io_in_stage(local_pes_7_11_io_in_stage),
    .io_out_q(local_pes_7_11_io_out_q),
    .io_out_sum(local_pes_7_11_io_out_sum),
    .io_out_sum_exp(local_pes_7_11_io_out_sum_exp),
    .io_out_kv(local_pes_7_11_io_out_kv),
    .io_out_stage(local_pes_7_11_io_out_stage)
  );
  PE_1 local_pes_7_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_12_clock),
    .reset(local_pes_7_12_reset),
    .io_in_q(local_pes_7_12_io_in_q),
    .io_in_sum(local_pes_7_12_io_in_sum),
    .io_in_sum_exp(local_pes_7_12_io_in_sum_exp),
    .io_in_kv(local_pes_7_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_12_io_in_inv_sum),
    .io_in_stage(local_pes_7_12_io_in_stage),
    .io_out_q(local_pes_7_12_io_out_q),
    .io_out_sum(local_pes_7_12_io_out_sum),
    .io_out_sum_exp(local_pes_7_12_io_out_sum_exp),
    .io_out_kv(local_pes_7_12_io_out_kv),
    .io_out_stage(local_pes_7_12_io_out_stage)
  );
  PE_1 local_pes_7_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_13_clock),
    .reset(local_pes_7_13_reset),
    .io_in_q(local_pes_7_13_io_in_q),
    .io_in_sum(local_pes_7_13_io_in_sum),
    .io_in_sum_exp(local_pes_7_13_io_in_sum_exp),
    .io_in_kv(local_pes_7_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_13_io_in_inv_sum),
    .io_in_stage(local_pes_7_13_io_in_stage),
    .io_out_q(local_pes_7_13_io_out_q),
    .io_out_sum(local_pes_7_13_io_out_sum),
    .io_out_sum_exp(local_pes_7_13_io_out_sum_exp),
    .io_out_kv(local_pes_7_13_io_out_kv),
    .io_out_stage(local_pes_7_13_io_out_stage)
  );
  PE_1 local_pes_7_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_14_clock),
    .reset(local_pes_7_14_reset),
    .io_in_q(local_pes_7_14_io_in_q),
    .io_in_sum(local_pes_7_14_io_in_sum),
    .io_in_sum_exp(local_pes_7_14_io_in_sum_exp),
    .io_in_kv(local_pes_7_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_14_io_in_inv_sum),
    .io_in_stage(local_pes_7_14_io_in_stage),
    .io_out_q(local_pes_7_14_io_out_q),
    .io_out_sum(local_pes_7_14_io_out_sum),
    .io_out_sum_exp(local_pes_7_14_io_out_sum_exp),
    .io_out_kv(local_pes_7_14_io_out_kv),
    .io_out_stage(local_pes_7_14_io_out_stage)
  );
  PE_1 local_pes_7_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_15_clock),
    .reset(local_pes_7_15_reset),
    .io_in_q(local_pes_7_15_io_in_q),
    .io_in_sum(local_pes_7_15_io_in_sum),
    .io_in_sum_exp(local_pes_7_15_io_in_sum_exp),
    .io_in_kv(local_pes_7_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_15_io_in_inv_sum),
    .io_in_stage(local_pes_7_15_io_in_stage),
    .io_out_q(local_pes_7_15_io_out_q),
    .io_out_sum(local_pes_7_15_io_out_sum),
    .io_out_sum_exp(local_pes_7_15_io_out_sum_exp),
    .io_out_kv(local_pes_7_15_io_out_kv),
    .io_out_stage(local_pes_7_15_io_out_stage)
  );
  PE_1 local_pes_7_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_16_clock),
    .reset(local_pes_7_16_reset),
    .io_in_q(local_pes_7_16_io_in_q),
    .io_in_sum(local_pes_7_16_io_in_sum),
    .io_in_sum_exp(local_pes_7_16_io_in_sum_exp),
    .io_in_kv(local_pes_7_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_16_io_in_inv_sum),
    .io_in_stage(local_pes_7_16_io_in_stage),
    .io_out_q(local_pes_7_16_io_out_q),
    .io_out_sum(local_pes_7_16_io_out_sum),
    .io_out_sum_exp(local_pes_7_16_io_out_sum_exp),
    .io_out_kv(local_pes_7_16_io_out_kv),
    .io_out_stage(local_pes_7_16_io_out_stage)
  );
  PE_1 local_pes_7_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_17_clock),
    .reset(local_pes_7_17_reset),
    .io_in_q(local_pes_7_17_io_in_q),
    .io_in_sum(local_pes_7_17_io_in_sum),
    .io_in_sum_exp(local_pes_7_17_io_in_sum_exp),
    .io_in_kv(local_pes_7_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_17_io_in_inv_sum),
    .io_in_stage(local_pes_7_17_io_in_stage),
    .io_out_q(local_pes_7_17_io_out_q),
    .io_out_sum(local_pes_7_17_io_out_sum),
    .io_out_sum_exp(local_pes_7_17_io_out_sum_exp),
    .io_out_kv(local_pes_7_17_io_out_kv),
    .io_out_stage(local_pes_7_17_io_out_stage)
  );
  PE_1 local_pes_7_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_18_clock),
    .reset(local_pes_7_18_reset),
    .io_in_q(local_pes_7_18_io_in_q),
    .io_in_sum(local_pes_7_18_io_in_sum),
    .io_in_sum_exp(local_pes_7_18_io_in_sum_exp),
    .io_in_kv(local_pes_7_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_18_io_in_inv_sum),
    .io_in_stage(local_pes_7_18_io_in_stage),
    .io_out_q(local_pes_7_18_io_out_q),
    .io_out_sum(local_pes_7_18_io_out_sum),
    .io_out_sum_exp(local_pes_7_18_io_out_sum_exp),
    .io_out_kv(local_pes_7_18_io_out_kv),
    .io_out_stage(local_pes_7_18_io_out_stage)
  );
  PE_1 local_pes_7_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_19_clock),
    .reset(local_pes_7_19_reset),
    .io_in_q(local_pes_7_19_io_in_q),
    .io_in_sum(local_pes_7_19_io_in_sum),
    .io_in_sum_exp(local_pes_7_19_io_in_sum_exp),
    .io_in_kv(local_pes_7_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_19_io_in_inv_sum),
    .io_in_stage(local_pes_7_19_io_in_stage),
    .io_out_q(local_pes_7_19_io_out_q),
    .io_out_sum(local_pes_7_19_io_out_sum),
    .io_out_sum_exp(local_pes_7_19_io_out_sum_exp),
    .io_out_kv(local_pes_7_19_io_out_kv),
    .io_out_stage(local_pes_7_19_io_out_stage)
  );
  PE_1 local_pes_7_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_20_clock),
    .reset(local_pes_7_20_reset),
    .io_in_q(local_pes_7_20_io_in_q),
    .io_in_sum(local_pes_7_20_io_in_sum),
    .io_in_sum_exp(local_pes_7_20_io_in_sum_exp),
    .io_in_kv(local_pes_7_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_20_io_in_inv_sum),
    .io_in_stage(local_pes_7_20_io_in_stage),
    .io_out_q(local_pes_7_20_io_out_q),
    .io_out_sum(local_pes_7_20_io_out_sum),
    .io_out_sum_exp(local_pes_7_20_io_out_sum_exp),
    .io_out_kv(local_pes_7_20_io_out_kv),
    .io_out_stage(local_pes_7_20_io_out_stage)
  );
  PE_1 local_pes_7_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_21_clock),
    .reset(local_pes_7_21_reset),
    .io_in_q(local_pes_7_21_io_in_q),
    .io_in_sum(local_pes_7_21_io_in_sum),
    .io_in_sum_exp(local_pes_7_21_io_in_sum_exp),
    .io_in_kv(local_pes_7_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_21_io_in_inv_sum),
    .io_in_stage(local_pes_7_21_io_in_stage),
    .io_out_q(local_pes_7_21_io_out_q),
    .io_out_sum(local_pes_7_21_io_out_sum),
    .io_out_sum_exp(local_pes_7_21_io_out_sum_exp),
    .io_out_kv(local_pes_7_21_io_out_kv),
    .io_out_stage(local_pes_7_21_io_out_stage)
  );
  PE_1 local_pes_7_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_22_clock),
    .reset(local_pes_7_22_reset),
    .io_in_q(local_pes_7_22_io_in_q),
    .io_in_sum(local_pes_7_22_io_in_sum),
    .io_in_sum_exp(local_pes_7_22_io_in_sum_exp),
    .io_in_kv(local_pes_7_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_22_io_in_inv_sum),
    .io_in_stage(local_pes_7_22_io_in_stage),
    .io_out_q(local_pes_7_22_io_out_q),
    .io_out_sum(local_pes_7_22_io_out_sum),
    .io_out_sum_exp(local_pes_7_22_io_out_sum_exp),
    .io_out_kv(local_pes_7_22_io_out_kv),
    .io_out_stage(local_pes_7_22_io_out_stage)
  );
  PE_1 local_pes_7_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_23_clock),
    .reset(local_pes_7_23_reset),
    .io_in_q(local_pes_7_23_io_in_q),
    .io_in_sum(local_pes_7_23_io_in_sum),
    .io_in_sum_exp(local_pes_7_23_io_in_sum_exp),
    .io_in_kv(local_pes_7_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_23_io_in_inv_sum),
    .io_in_stage(local_pes_7_23_io_in_stage),
    .io_out_q(local_pes_7_23_io_out_q),
    .io_out_sum(local_pes_7_23_io_out_sum),
    .io_out_sum_exp(local_pes_7_23_io_out_sum_exp),
    .io_out_kv(local_pes_7_23_io_out_kv),
    .io_out_stage(local_pes_7_23_io_out_stage)
  );
  PE_1 local_pes_7_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_24_clock),
    .reset(local_pes_7_24_reset),
    .io_in_q(local_pes_7_24_io_in_q),
    .io_in_sum(local_pes_7_24_io_in_sum),
    .io_in_sum_exp(local_pes_7_24_io_in_sum_exp),
    .io_in_kv(local_pes_7_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_24_io_in_inv_sum),
    .io_in_stage(local_pes_7_24_io_in_stage),
    .io_out_q(local_pes_7_24_io_out_q),
    .io_out_sum(local_pes_7_24_io_out_sum),
    .io_out_sum_exp(local_pes_7_24_io_out_sum_exp),
    .io_out_kv(local_pes_7_24_io_out_kv),
    .io_out_stage(local_pes_7_24_io_out_stage)
  );
  PE_1 local_pes_7_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_25_clock),
    .reset(local_pes_7_25_reset),
    .io_in_q(local_pes_7_25_io_in_q),
    .io_in_sum(local_pes_7_25_io_in_sum),
    .io_in_sum_exp(local_pes_7_25_io_in_sum_exp),
    .io_in_kv(local_pes_7_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_25_io_in_inv_sum),
    .io_in_stage(local_pes_7_25_io_in_stage),
    .io_out_q(local_pes_7_25_io_out_q),
    .io_out_sum(local_pes_7_25_io_out_sum),
    .io_out_sum_exp(local_pes_7_25_io_out_sum_exp),
    .io_out_kv(local_pes_7_25_io_out_kv),
    .io_out_stage(local_pes_7_25_io_out_stage)
  );
  PE_1 local_pes_7_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_26_clock),
    .reset(local_pes_7_26_reset),
    .io_in_q(local_pes_7_26_io_in_q),
    .io_in_sum(local_pes_7_26_io_in_sum),
    .io_in_sum_exp(local_pes_7_26_io_in_sum_exp),
    .io_in_kv(local_pes_7_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_26_io_in_inv_sum),
    .io_in_stage(local_pes_7_26_io_in_stage),
    .io_out_q(local_pes_7_26_io_out_q),
    .io_out_sum(local_pes_7_26_io_out_sum),
    .io_out_sum_exp(local_pes_7_26_io_out_sum_exp),
    .io_out_kv(local_pes_7_26_io_out_kv),
    .io_out_stage(local_pes_7_26_io_out_stage)
  );
  PE_1 local_pes_7_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_27_clock),
    .reset(local_pes_7_27_reset),
    .io_in_q(local_pes_7_27_io_in_q),
    .io_in_sum(local_pes_7_27_io_in_sum),
    .io_in_sum_exp(local_pes_7_27_io_in_sum_exp),
    .io_in_kv(local_pes_7_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_27_io_in_inv_sum),
    .io_in_stage(local_pes_7_27_io_in_stage),
    .io_out_q(local_pes_7_27_io_out_q),
    .io_out_sum(local_pes_7_27_io_out_sum),
    .io_out_sum_exp(local_pes_7_27_io_out_sum_exp),
    .io_out_kv(local_pes_7_27_io_out_kv),
    .io_out_stage(local_pes_7_27_io_out_stage)
  );
  PE_1 local_pes_7_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_28_clock),
    .reset(local_pes_7_28_reset),
    .io_in_q(local_pes_7_28_io_in_q),
    .io_in_sum(local_pes_7_28_io_in_sum),
    .io_in_sum_exp(local_pes_7_28_io_in_sum_exp),
    .io_in_kv(local_pes_7_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_28_io_in_inv_sum),
    .io_in_stage(local_pes_7_28_io_in_stage),
    .io_out_q(local_pes_7_28_io_out_q),
    .io_out_sum(local_pes_7_28_io_out_sum),
    .io_out_sum_exp(local_pes_7_28_io_out_sum_exp),
    .io_out_kv(local_pes_7_28_io_out_kv),
    .io_out_stage(local_pes_7_28_io_out_stage)
  );
  PE_1 local_pes_7_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_29_clock),
    .reset(local_pes_7_29_reset),
    .io_in_q(local_pes_7_29_io_in_q),
    .io_in_sum(local_pes_7_29_io_in_sum),
    .io_in_sum_exp(local_pes_7_29_io_in_sum_exp),
    .io_in_kv(local_pes_7_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_29_io_in_inv_sum),
    .io_in_stage(local_pes_7_29_io_in_stage),
    .io_out_q(local_pes_7_29_io_out_q),
    .io_out_sum(local_pes_7_29_io_out_sum),
    .io_out_sum_exp(local_pes_7_29_io_out_sum_exp),
    .io_out_kv(local_pes_7_29_io_out_kv),
    .io_out_stage(local_pes_7_29_io_out_stage)
  );
  PE_1 local_pes_7_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_30_clock),
    .reset(local_pes_7_30_reset),
    .io_in_q(local_pes_7_30_io_in_q),
    .io_in_sum(local_pes_7_30_io_in_sum),
    .io_in_sum_exp(local_pes_7_30_io_in_sum_exp),
    .io_in_kv(local_pes_7_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_30_io_in_inv_sum),
    .io_in_stage(local_pes_7_30_io_in_stage),
    .io_out_q(local_pes_7_30_io_out_q),
    .io_out_sum(local_pes_7_30_io_out_sum),
    .io_out_sum_exp(local_pes_7_30_io_out_sum_exp),
    .io_out_kv(local_pes_7_30_io_out_kv),
    .io_out_stage(local_pes_7_30_io_out_stage)
  );
  PE_1 local_pes_7_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_7_31_clock),
    .reset(local_pes_7_31_reset),
    .io_in_q(local_pes_7_31_io_in_q),
    .io_in_sum(local_pes_7_31_io_in_sum),
    .io_in_sum_exp(local_pes_7_31_io_in_sum_exp),
    .io_in_kv(local_pes_7_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_7_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_7_31_io_in_inv_sum),
    .io_in_stage(local_pes_7_31_io_in_stage),
    .io_out_q(local_pes_7_31_io_out_q),
    .io_out_sum(local_pes_7_31_io_out_sum),
    .io_out_sum_exp(local_pes_7_31_io_out_sum_exp),
    .io_out_kv(local_pes_7_31_io_out_kv),
    .io_out_stage(local_pes_7_31_io_out_stage)
  );
  PE local_pes_8_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_0_clock),
    .reset(local_pes_8_0_reset),
    .io_in_q(local_pes_8_0_io_in_q),
    .io_in_kv(local_pes_8_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_0_io_in_inv_sum),
    .io_in_stage(local_pes_8_0_io_in_stage),
    .io_out_q(local_pes_8_0_io_out_q),
    .io_out_sum(local_pes_8_0_io_out_sum),
    .io_out_kv(local_pes_8_0_io_out_kv),
    .io_out_stage(local_pes_8_0_io_out_stage)
  );
  PE_1 local_pes_8_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_1_clock),
    .reset(local_pes_8_1_reset),
    .io_in_q(local_pes_8_1_io_in_q),
    .io_in_sum(local_pes_8_1_io_in_sum),
    .io_in_sum_exp(local_pes_8_1_io_in_sum_exp),
    .io_in_kv(local_pes_8_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_1_io_in_inv_sum),
    .io_in_stage(local_pes_8_1_io_in_stage),
    .io_out_q(local_pes_8_1_io_out_q),
    .io_out_sum(local_pes_8_1_io_out_sum),
    .io_out_sum_exp(local_pes_8_1_io_out_sum_exp),
    .io_out_kv(local_pes_8_1_io_out_kv),
    .io_out_stage(local_pes_8_1_io_out_stage)
  );
  PE_1 local_pes_8_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_2_clock),
    .reset(local_pes_8_2_reset),
    .io_in_q(local_pes_8_2_io_in_q),
    .io_in_sum(local_pes_8_2_io_in_sum),
    .io_in_sum_exp(local_pes_8_2_io_in_sum_exp),
    .io_in_kv(local_pes_8_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_2_io_in_inv_sum),
    .io_in_stage(local_pes_8_2_io_in_stage),
    .io_out_q(local_pes_8_2_io_out_q),
    .io_out_sum(local_pes_8_2_io_out_sum),
    .io_out_sum_exp(local_pes_8_2_io_out_sum_exp),
    .io_out_kv(local_pes_8_2_io_out_kv),
    .io_out_stage(local_pes_8_2_io_out_stage)
  );
  PE_1 local_pes_8_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_3_clock),
    .reset(local_pes_8_3_reset),
    .io_in_q(local_pes_8_3_io_in_q),
    .io_in_sum(local_pes_8_3_io_in_sum),
    .io_in_sum_exp(local_pes_8_3_io_in_sum_exp),
    .io_in_kv(local_pes_8_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_3_io_in_inv_sum),
    .io_in_stage(local_pes_8_3_io_in_stage),
    .io_out_q(local_pes_8_3_io_out_q),
    .io_out_sum(local_pes_8_3_io_out_sum),
    .io_out_sum_exp(local_pes_8_3_io_out_sum_exp),
    .io_out_kv(local_pes_8_3_io_out_kv),
    .io_out_stage(local_pes_8_3_io_out_stage)
  );
  PE_1 local_pes_8_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_4_clock),
    .reset(local_pes_8_4_reset),
    .io_in_q(local_pes_8_4_io_in_q),
    .io_in_sum(local_pes_8_4_io_in_sum),
    .io_in_sum_exp(local_pes_8_4_io_in_sum_exp),
    .io_in_kv(local_pes_8_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_4_io_in_inv_sum),
    .io_in_stage(local_pes_8_4_io_in_stage),
    .io_out_q(local_pes_8_4_io_out_q),
    .io_out_sum(local_pes_8_4_io_out_sum),
    .io_out_sum_exp(local_pes_8_4_io_out_sum_exp),
    .io_out_kv(local_pes_8_4_io_out_kv),
    .io_out_stage(local_pes_8_4_io_out_stage)
  );
  PE_1 local_pes_8_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_5_clock),
    .reset(local_pes_8_5_reset),
    .io_in_q(local_pes_8_5_io_in_q),
    .io_in_sum(local_pes_8_5_io_in_sum),
    .io_in_sum_exp(local_pes_8_5_io_in_sum_exp),
    .io_in_kv(local_pes_8_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_5_io_in_inv_sum),
    .io_in_stage(local_pes_8_5_io_in_stage),
    .io_out_q(local_pes_8_5_io_out_q),
    .io_out_sum(local_pes_8_5_io_out_sum),
    .io_out_sum_exp(local_pes_8_5_io_out_sum_exp),
    .io_out_kv(local_pes_8_5_io_out_kv),
    .io_out_stage(local_pes_8_5_io_out_stage)
  );
  PE_1 local_pes_8_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_6_clock),
    .reset(local_pes_8_6_reset),
    .io_in_q(local_pes_8_6_io_in_q),
    .io_in_sum(local_pes_8_6_io_in_sum),
    .io_in_sum_exp(local_pes_8_6_io_in_sum_exp),
    .io_in_kv(local_pes_8_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_6_io_in_inv_sum),
    .io_in_stage(local_pes_8_6_io_in_stage),
    .io_out_q(local_pes_8_6_io_out_q),
    .io_out_sum(local_pes_8_6_io_out_sum),
    .io_out_sum_exp(local_pes_8_6_io_out_sum_exp),
    .io_out_kv(local_pes_8_6_io_out_kv),
    .io_out_stage(local_pes_8_6_io_out_stage)
  );
  PE_1 local_pes_8_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_7_clock),
    .reset(local_pes_8_7_reset),
    .io_in_q(local_pes_8_7_io_in_q),
    .io_in_sum(local_pes_8_7_io_in_sum),
    .io_in_sum_exp(local_pes_8_7_io_in_sum_exp),
    .io_in_kv(local_pes_8_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_7_io_in_inv_sum),
    .io_in_stage(local_pes_8_7_io_in_stage),
    .io_out_q(local_pes_8_7_io_out_q),
    .io_out_sum(local_pes_8_7_io_out_sum),
    .io_out_sum_exp(local_pes_8_7_io_out_sum_exp),
    .io_out_kv(local_pes_8_7_io_out_kv),
    .io_out_stage(local_pes_8_7_io_out_stage)
  );
  PE_1 local_pes_8_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_8_clock),
    .reset(local_pes_8_8_reset),
    .io_in_q(local_pes_8_8_io_in_q),
    .io_in_sum(local_pes_8_8_io_in_sum),
    .io_in_sum_exp(local_pes_8_8_io_in_sum_exp),
    .io_in_kv(local_pes_8_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_8_io_in_inv_sum),
    .io_in_stage(local_pes_8_8_io_in_stage),
    .io_out_q(local_pes_8_8_io_out_q),
    .io_out_sum(local_pes_8_8_io_out_sum),
    .io_out_sum_exp(local_pes_8_8_io_out_sum_exp),
    .io_out_kv(local_pes_8_8_io_out_kv),
    .io_out_stage(local_pes_8_8_io_out_stage)
  );
  PE_1 local_pes_8_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_9_clock),
    .reset(local_pes_8_9_reset),
    .io_in_q(local_pes_8_9_io_in_q),
    .io_in_sum(local_pes_8_9_io_in_sum),
    .io_in_sum_exp(local_pes_8_9_io_in_sum_exp),
    .io_in_kv(local_pes_8_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_9_io_in_inv_sum),
    .io_in_stage(local_pes_8_9_io_in_stage),
    .io_out_q(local_pes_8_9_io_out_q),
    .io_out_sum(local_pes_8_9_io_out_sum),
    .io_out_sum_exp(local_pes_8_9_io_out_sum_exp),
    .io_out_kv(local_pes_8_9_io_out_kv),
    .io_out_stage(local_pes_8_9_io_out_stage)
  );
  PE_1 local_pes_8_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_10_clock),
    .reset(local_pes_8_10_reset),
    .io_in_q(local_pes_8_10_io_in_q),
    .io_in_sum(local_pes_8_10_io_in_sum),
    .io_in_sum_exp(local_pes_8_10_io_in_sum_exp),
    .io_in_kv(local_pes_8_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_10_io_in_inv_sum),
    .io_in_stage(local_pes_8_10_io_in_stage),
    .io_out_q(local_pes_8_10_io_out_q),
    .io_out_sum(local_pes_8_10_io_out_sum),
    .io_out_sum_exp(local_pes_8_10_io_out_sum_exp),
    .io_out_kv(local_pes_8_10_io_out_kv),
    .io_out_stage(local_pes_8_10_io_out_stage)
  );
  PE_1 local_pes_8_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_11_clock),
    .reset(local_pes_8_11_reset),
    .io_in_q(local_pes_8_11_io_in_q),
    .io_in_sum(local_pes_8_11_io_in_sum),
    .io_in_sum_exp(local_pes_8_11_io_in_sum_exp),
    .io_in_kv(local_pes_8_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_11_io_in_inv_sum),
    .io_in_stage(local_pes_8_11_io_in_stage),
    .io_out_q(local_pes_8_11_io_out_q),
    .io_out_sum(local_pes_8_11_io_out_sum),
    .io_out_sum_exp(local_pes_8_11_io_out_sum_exp),
    .io_out_kv(local_pes_8_11_io_out_kv),
    .io_out_stage(local_pes_8_11_io_out_stage)
  );
  PE_1 local_pes_8_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_12_clock),
    .reset(local_pes_8_12_reset),
    .io_in_q(local_pes_8_12_io_in_q),
    .io_in_sum(local_pes_8_12_io_in_sum),
    .io_in_sum_exp(local_pes_8_12_io_in_sum_exp),
    .io_in_kv(local_pes_8_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_12_io_in_inv_sum),
    .io_in_stage(local_pes_8_12_io_in_stage),
    .io_out_q(local_pes_8_12_io_out_q),
    .io_out_sum(local_pes_8_12_io_out_sum),
    .io_out_sum_exp(local_pes_8_12_io_out_sum_exp),
    .io_out_kv(local_pes_8_12_io_out_kv),
    .io_out_stage(local_pes_8_12_io_out_stage)
  );
  PE_1 local_pes_8_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_13_clock),
    .reset(local_pes_8_13_reset),
    .io_in_q(local_pes_8_13_io_in_q),
    .io_in_sum(local_pes_8_13_io_in_sum),
    .io_in_sum_exp(local_pes_8_13_io_in_sum_exp),
    .io_in_kv(local_pes_8_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_13_io_in_inv_sum),
    .io_in_stage(local_pes_8_13_io_in_stage),
    .io_out_q(local_pes_8_13_io_out_q),
    .io_out_sum(local_pes_8_13_io_out_sum),
    .io_out_sum_exp(local_pes_8_13_io_out_sum_exp),
    .io_out_kv(local_pes_8_13_io_out_kv),
    .io_out_stage(local_pes_8_13_io_out_stage)
  );
  PE_1 local_pes_8_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_14_clock),
    .reset(local_pes_8_14_reset),
    .io_in_q(local_pes_8_14_io_in_q),
    .io_in_sum(local_pes_8_14_io_in_sum),
    .io_in_sum_exp(local_pes_8_14_io_in_sum_exp),
    .io_in_kv(local_pes_8_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_14_io_in_inv_sum),
    .io_in_stage(local_pes_8_14_io_in_stage),
    .io_out_q(local_pes_8_14_io_out_q),
    .io_out_sum(local_pes_8_14_io_out_sum),
    .io_out_sum_exp(local_pes_8_14_io_out_sum_exp),
    .io_out_kv(local_pes_8_14_io_out_kv),
    .io_out_stage(local_pes_8_14_io_out_stage)
  );
  PE_1 local_pes_8_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_15_clock),
    .reset(local_pes_8_15_reset),
    .io_in_q(local_pes_8_15_io_in_q),
    .io_in_sum(local_pes_8_15_io_in_sum),
    .io_in_sum_exp(local_pes_8_15_io_in_sum_exp),
    .io_in_kv(local_pes_8_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_15_io_in_inv_sum),
    .io_in_stage(local_pes_8_15_io_in_stage),
    .io_out_q(local_pes_8_15_io_out_q),
    .io_out_sum(local_pes_8_15_io_out_sum),
    .io_out_sum_exp(local_pes_8_15_io_out_sum_exp),
    .io_out_kv(local_pes_8_15_io_out_kv),
    .io_out_stage(local_pes_8_15_io_out_stage)
  );
  PE_1 local_pes_8_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_16_clock),
    .reset(local_pes_8_16_reset),
    .io_in_q(local_pes_8_16_io_in_q),
    .io_in_sum(local_pes_8_16_io_in_sum),
    .io_in_sum_exp(local_pes_8_16_io_in_sum_exp),
    .io_in_kv(local_pes_8_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_16_io_in_inv_sum),
    .io_in_stage(local_pes_8_16_io_in_stage),
    .io_out_q(local_pes_8_16_io_out_q),
    .io_out_sum(local_pes_8_16_io_out_sum),
    .io_out_sum_exp(local_pes_8_16_io_out_sum_exp),
    .io_out_kv(local_pes_8_16_io_out_kv),
    .io_out_stage(local_pes_8_16_io_out_stage)
  );
  PE_1 local_pes_8_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_17_clock),
    .reset(local_pes_8_17_reset),
    .io_in_q(local_pes_8_17_io_in_q),
    .io_in_sum(local_pes_8_17_io_in_sum),
    .io_in_sum_exp(local_pes_8_17_io_in_sum_exp),
    .io_in_kv(local_pes_8_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_17_io_in_inv_sum),
    .io_in_stage(local_pes_8_17_io_in_stage),
    .io_out_q(local_pes_8_17_io_out_q),
    .io_out_sum(local_pes_8_17_io_out_sum),
    .io_out_sum_exp(local_pes_8_17_io_out_sum_exp),
    .io_out_kv(local_pes_8_17_io_out_kv),
    .io_out_stage(local_pes_8_17_io_out_stage)
  );
  PE_1 local_pes_8_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_18_clock),
    .reset(local_pes_8_18_reset),
    .io_in_q(local_pes_8_18_io_in_q),
    .io_in_sum(local_pes_8_18_io_in_sum),
    .io_in_sum_exp(local_pes_8_18_io_in_sum_exp),
    .io_in_kv(local_pes_8_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_18_io_in_inv_sum),
    .io_in_stage(local_pes_8_18_io_in_stage),
    .io_out_q(local_pes_8_18_io_out_q),
    .io_out_sum(local_pes_8_18_io_out_sum),
    .io_out_sum_exp(local_pes_8_18_io_out_sum_exp),
    .io_out_kv(local_pes_8_18_io_out_kv),
    .io_out_stage(local_pes_8_18_io_out_stage)
  );
  PE_1 local_pes_8_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_19_clock),
    .reset(local_pes_8_19_reset),
    .io_in_q(local_pes_8_19_io_in_q),
    .io_in_sum(local_pes_8_19_io_in_sum),
    .io_in_sum_exp(local_pes_8_19_io_in_sum_exp),
    .io_in_kv(local_pes_8_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_19_io_in_inv_sum),
    .io_in_stage(local_pes_8_19_io_in_stage),
    .io_out_q(local_pes_8_19_io_out_q),
    .io_out_sum(local_pes_8_19_io_out_sum),
    .io_out_sum_exp(local_pes_8_19_io_out_sum_exp),
    .io_out_kv(local_pes_8_19_io_out_kv),
    .io_out_stage(local_pes_8_19_io_out_stage)
  );
  PE_1 local_pes_8_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_20_clock),
    .reset(local_pes_8_20_reset),
    .io_in_q(local_pes_8_20_io_in_q),
    .io_in_sum(local_pes_8_20_io_in_sum),
    .io_in_sum_exp(local_pes_8_20_io_in_sum_exp),
    .io_in_kv(local_pes_8_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_20_io_in_inv_sum),
    .io_in_stage(local_pes_8_20_io_in_stage),
    .io_out_q(local_pes_8_20_io_out_q),
    .io_out_sum(local_pes_8_20_io_out_sum),
    .io_out_sum_exp(local_pes_8_20_io_out_sum_exp),
    .io_out_kv(local_pes_8_20_io_out_kv),
    .io_out_stage(local_pes_8_20_io_out_stage)
  );
  PE_1 local_pes_8_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_21_clock),
    .reset(local_pes_8_21_reset),
    .io_in_q(local_pes_8_21_io_in_q),
    .io_in_sum(local_pes_8_21_io_in_sum),
    .io_in_sum_exp(local_pes_8_21_io_in_sum_exp),
    .io_in_kv(local_pes_8_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_21_io_in_inv_sum),
    .io_in_stage(local_pes_8_21_io_in_stage),
    .io_out_q(local_pes_8_21_io_out_q),
    .io_out_sum(local_pes_8_21_io_out_sum),
    .io_out_sum_exp(local_pes_8_21_io_out_sum_exp),
    .io_out_kv(local_pes_8_21_io_out_kv),
    .io_out_stage(local_pes_8_21_io_out_stage)
  );
  PE_1 local_pes_8_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_22_clock),
    .reset(local_pes_8_22_reset),
    .io_in_q(local_pes_8_22_io_in_q),
    .io_in_sum(local_pes_8_22_io_in_sum),
    .io_in_sum_exp(local_pes_8_22_io_in_sum_exp),
    .io_in_kv(local_pes_8_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_22_io_in_inv_sum),
    .io_in_stage(local_pes_8_22_io_in_stage),
    .io_out_q(local_pes_8_22_io_out_q),
    .io_out_sum(local_pes_8_22_io_out_sum),
    .io_out_sum_exp(local_pes_8_22_io_out_sum_exp),
    .io_out_kv(local_pes_8_22_io_out_kv),
    .io_out_stage(local_pes_8_22_io_out_stage)
  );
  PE_1 local_pes_8_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_23_clock),
    .reset(local_pes_8_23_reset),
    .io_in_q(local_pes_8_23_io_in_q),
    .io_in_sum(local_pes_8_23_io_in_sum),
    .io_in_sum_exp(local_pes_8_23_io_in_sum_exp),
    .io_in_kv(local_pes_8_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_23_io_in_inv_sum),
    .io_in_stage(local_pes_8_23_io_in_stage),
    .io_out_q(local_pes_8_23_io_out_q),
    .io_out_sum(local_pes_8_23_io_out_sum),
    .io_out_sum_exp(local_pes_8_23_io_out_sum_exp),
    .io_out_kv(local_pes_8_23_io_out_kv),
    .io_out_stage(local_pes_8_23_io_out_stage)
  );
  PE_1 local_pes_8_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_24_clock),
    .reset(local_pes_8_24_reset),
    .io_in_q(local_pes_8_24_io_in_q),
    .io_in_sum(local_pes_8_24_io_in_sum),
    .io_in_sum_exp(local_pes_8_24_io_in_sum_exp),
    .io_in_kv(local_pes_8_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_24_io_in_inv_sum),
    .io_in_stage(local_pes_8_24_io_in_stage),
    .io_out_q(local_pes_8_24_io_out_q),
    .io_out_sum(local_pes_8_24_io_out_sum),
    .io_out_sum_exp(local_pes_8_24_io_out_sum_exp),
    .io_out_kv(local_pes_8_24_io_out_kv),
    .io_out_stage(local_pes_8_24_io_out_stage)
  );
  PE_1 local_pes_8_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_25_clock),
    .reset(local_pes_8_25_reset),
    .io_in_q(local_pes_8_25_io_in_q),
    .io_in_sum(local_pes_8_25_io_in_sum),
    .io_in_sum_exp(local_pes_8_25_io_in_sum_exp),
    .io_in_kv(local_pes_8_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_25_io_in_inv_sum),
    .io_in_stage(local_pes_8_25_io_in_stage),
    .io_out_q(local_pes_8_25_io_out_q),
    .io_out_sum(local_pes_8_25_io_out_sum),
    .io_out_sum_exp(local_pes_8_25_io_out_sum_exp),
    .io_out_kv(local_pes_8_25_io_out_kv),
    .io_out_stage(local_pes_8_25_io_out_stage)
  );
  PE_1 local_pes_8_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_26_clock),
    .reset(local_pes_8_26_reset),
    .io_in_q(local_pes_8_26_io_in_q),
    .io_in_sum(local_pes_8_26_io_in_sum),
    .io_in_sum_exp(local_pes_8_26_io_in_sum_exp),
    .io_in_kv(local_pes_8_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_26_io_in_inv_sum),
    .io_in_stage(local_pes_8_26_io_in_stage),
    .io_out_q(local_pes_8_26_io_out_q),
    .io_out_sum(local_pes_8_26_io_out_sum),
    .io_out_sum_exp(local_pes_8_26_io_out_sum_exp),
    .io_out_kv(local_pes_8_26_io_out_kv),
    .io_out_stage(local_pes_8_26_io_out_stage)
  );
  PE_1 local_pes_8_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_27_clock),
    .reset(local_pes_8_27_reset),
    .io_in_q(local_pes_8_27_io_in_q),
    .io_in_sum(local_pes_8_27_io_in_sum),
    .io_in_sum_exp(local_pes_8_27_io_in_sum_exp),
    .io_in_kv(local_pes_8_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_27_io_in_inv_sum),
    .io_in_stage(local_pes_8_27_io_in_stage),
    .io_out_q(local_pes_8_27_io_out_q),
    .io_out_sum(local_pes_8_27_io_out_sum),
    .io_out_sum_exp(local_pes_8_27_io_out_sum_exp),
    .io_out_kv(local_pes_8_27_io_out_kv),
    .io_out_stage(local_pes_8_27_io_out_stage)
  );
  PE_1 local_pes_8_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_28_clock),
    .reset(local_pes_8_28_reset),
    .io_in_q(local_pes_8_28_io_in_q),
    .io_in_sum(local_pes_8_28_io_in_sum),
    .io_in_sum_exp(local_pes_8_28_io_in_sum_exp),
    .io_in_kv(local_pes_8_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_28_io_in_inv_sum),
    .io_in_stage(local_pes_8_28_io_in_stage),
    .io_out_q(local_pes_8_28_io_out_q),
    .io_out_sum(local_pes_8_28_io_out_sum),
    .io_out_sum_exp(local_pes_8_28_io_out_sum_exp),
    .io_out_kv(local_pes_8_28_io_out_kv),
    .io_out_stage(local_pes_8_28_io_out_stage)
  );
  PE_1 local_pes_8_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_29_clock),
    .reset(local_pes_8_29_reset),
    .io_in_q(local_pes_8_29_io_in_q),
    .io_in_sum(local_pes_8_29_io_in_sum),
    .io_in_sum_exp(local_pes_8_29_io_in_sum_exp),
    .io_in_kv(local_pes_8_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_29_io_in_inv_sum),
    .io_in_stage(local_pes_8_29_io_in_stage),
    .io_out_q(local_pes_8_29_io_out_q),
    .io_out_sum(local_pes_8_29_io_out_sum),
    .io_out_sum_exp(local_pes_8_29_io_out_sum_exp),
    .io_out_kv(local_pes_8_29_io_out_kv),
    .io_out_stage(local_pes_8_29_io_out_stage)
  );
  PE_1 local_pes_8_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_30_clock),
    .reset(local_pes_8_30_reset),
    .io_in_q(local_pes_8_30_io_in_q),
    .io_in_sum(local_pes_8_30_io_in_sum),
    .io_in_sum_exp(local_pes_8_30_io_in_sum_exp),
    .io_in_kv(local_pes_8_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_30_io_in_inv_sum),
    .io_in_stage(local_pes_8_30_io_in_stage),
    .io_out_q(local_pes_8_30_io_out_q),
    .io_out_sum(local_pes_8_30_io_out_sum),
    .io_out_sum_exp(local_pes_8_30_io_out_sum_exp),
    .io_out_kv(local_pes_8_30_io_out_kv),
    .io_out_stage(local_pes_8_30_io_out_stage)
  );
  PE_1 local_pes_8_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_8_31_clock),
    .reset(local_pes_8_31_reset),
    .io_in_q(local_pes_8_31_io_in_q),
    .io_in_sum(local_pes_8_31_io_in_sum),
    .io_in_sum_exp(local_pes_8_31_io_in_sum_exp),
    .io_in_kv(local_pes_8_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_8_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_8_31_io_in_inv_sum),
    .io_in_stage(local_pes_8_31_io_in_stage),
    .io_out_q(local_pes_8_31_io_out_q),
    .io_out_sum(local_pes_8_31_io_out_sum),
    .io_out_sum_exp(local_pes_8_31_io_out_sum_exp),
    .io_out_kv(local_pes_8_31_io_out_kv),
    .io_out_stage(local_pes_8_31_io_out_stage)
  );
  PE local_pes_9_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_0_clock),
    .reset(local_pes_9_0_reset),
    .io_in_q(local_pes_9_0_io_in_q),
    .io_in_kv(local_pes_9_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_0_io_in_inv_sum),
    .io_in_stage(local_pes_9_0_io_in_stage),
    .io_out_q(local_pes_9_0_io_out_q),
    .io_out_sum(local_pes_9_0_io_out_sum),
    .io_out_kv(local_pes_9_0_io_out_kv),
    .io_out_stage(local_pes_9_0_io_out_stage)
  );
  PE_1 local_pes_9_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_1_clock),
    .reset(local_pes_9_1_reset),
    .io_in_q(local_pes_9_1_io_in_q),
    .io_in_sum(local_pes_9_1_io_in_sum),
    .io_in_sum_exp(local_pes_9_1_io_in_sum_exp),
    .io_in_kv(local_pes_9_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_1_io_in_inv_sum),
    .io_in_stage(local_pes_9_1_io_in_stage),
    .io_out_q(local_pes_9_1_io_out_q),
    .io_out_sum(local_pes_9_1_io_out_sum),
    .io_out_sum_exp(local_pes_9_1_io_out_sum_exp),
    .io_out_kv(local_pes_9_1_io_out_kv),
    .io_out_stage(local_pes_9_1_io_out_stage)
  );
  PE_1 local_pes_9_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_2_clock),
    .reset(local_pes_9_2_reset),
    .io_in_q(local_pes_9_2_io_in_q),
    .io_in_sum(local_pes_9_2_io_in_sum),
    .io_in_sum_exp(local_pes_9_2_io_in_sum_exp),
    .io_in_kv(local_pes_9_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_2_io_in_inv_sum),
    .io_in_stage(local_pes_9_2_io_in_stage),
    .io_out_q(local_pes_9_2_io_out_q),
    .io_out_sum(local_pes_9_2_io_out_sum),
    .io_out_sum_exp(local_pes_9_2_io_out_sum_exp),
    .io_out_kv(local_pes_9_2_io_out_kv),
    .io_out_stage(local_pes_9_2_io_out_stage)
  );
  PE_1 local_pes_9_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_3_clock),
    .reset(local_pes_9_3_reset),
    .io_in_q(local_pes_9_3_io_in_q),
    .io_in_sum(local_pes_9_3_io_in_sum),
    .io_in_sum_exp(local_pes_9_3_io_in_sum_exp),
    .io_in_kv(local_pes_9_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_3_io_in_inv_sum),
    .io_in_stage(local_pes_9_3_io_in_stage),
    .io_out_q(local_pes_9_3_io_out_q),
    .io_out_sum(local_pes_9_3_io_out_sum),
    .io_out_sum_exp(local_pes_9_3_io_out_sum_exp),
    .io_out_kv(local_pes_9_3_io_out_kv),
    .io_out_stage(local_pes_9_3_io_out_stage)
  );
  PE_1 local_pes_9_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_4_clock),
    .reset(local_pes_9_4_reset),
    .io_in_q(local_pes_9_4_io_in_q),
    .io_in_sum(local_pes_9_4_io_in_sum),
    .io_in_sum_exp(local_pes_9_4_io_in_sum_exp),
    .io_in_kv(local_pes_9_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_4_io_in_inv_sum),
    .io_in_stage(local_pes_9_4_io_in_stage),
    .io_out_q(local_pes_9_4_io_out_q),
    .io_out_sum(local_pes_9_4_io_out_sum),
    .io_out_sum_exp(local_pes_9_4_io_out_sum_exp),
    .io_out_kv(local_pes_9_4_io_out_kv),
    .io_out_stage(local_pes_9_4_io_out_stage)
  );
  PE_1 local_pes_9_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_5_clock),
    .reset(local_pes_9_5_reset),
    .io_in_q(local_pes_9_5_io_in_q),
    .io_in_sum(local_pes_9_5_io_in_sum),
    .io_in_sum_exp(local_pes_9_5_io_in_sum_exp),
    .io_in_kv(local_pes_9_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_5_io_in_inv_sum),
    .io_in_stage(local_pes_9_5_io_in_stage),
    .io_out_q(local_pes_9_5_io_out_q),
    .io_out_sum(local_pes_9_5_io_out_sum),
    .io_out_sum_exp(local_pes_9_5_io_out_sum_exp),
    .io_out_kv(local_pes_9_5_io_out_kv),
    .io_out_stage(local_pes_9_5_io_out_stage)
  );
  PE_1 local_pes_9_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_6_clock),
    .reset(local_pes_9_6_reset),
    .io_in_q(local_pes_9_6_io_in_q),
    .io_in_sum(local_pes_9_6_io_in_sum),
    .io_in_sum_exp(local_pes_9_6_io_in_sum_exp),
    .io_in_kv(local_pes_9_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_6_io_in_inv_sum),
    .io_in_stage(local_pes_9_6_io_in_stage),
    .io_out_q(local_pes_9_6_io_out_q),
    .io_out_sum(local_pes_9_6_io_out_sum),
    .io_out_sum_exp(local_pes_9_6_io_out_sum_exp),
    .io_out_kv(local_pes_9_6_io_out_kv),
    .io_out_stage(local_pes_9_6_io_out_stage)
  );
  PE_1 local_pes_9_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_7_clock),
    .reset(local_pes_9_7_reset),
    .io_in_q(local_pes_9_7_io_in_q),
    .io_in_sum(local_pes_9_7_io_in_sum),
    .io_in_sum_exp(local_pes_9_7_io_in_sum_exp),
    .io_in_kv(local_pes_9_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_7_io_in_inv_sum),
    .io_in_stage(local_pes_9_7_io_in_stage),
    .io_out_q(local_pes_9_7_io_out_q),
    .io_out_sum(local_pes_9_7_io_out_sum),
    .io_out_sum_exp(local_pes_9_7_io_out_sum_exp),
    .io_out_kv(local_pes_9_7_io_out_kv),
    .io_out_stage(local_pes_9_7_io_out_stage)
  );
  PE_1 local_pes_9_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_8_clock),
    .reset(local_pes_9_8_reset),
    .io_in_q(local_pes_9_8_io_in_q),
    .io_in_sum(local_pes_9_8_io_in_sum),
    .io_in_sum_exp(local_pes_9_8_io_in_sum_exp),
    .io_in_kv(local_pes_9_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_8_io_in_inv_sum),
    .io_in_stage(local_pes_9_8_io_in_stage),
    .io_out_q(local_pes_9_8_io_out_q),
    .io_out_sum(local_pes_9_8_io_out_sum),
    .io_out_sum_exp(local_pes_9_8_io_out_sum_exp),
    .io_out_kv(local_pes_9_8_io_out_kv),
    .io_out_stage(local_pes_9_8_io_out_stage)
  );
  PE_1 local_pes_9_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_9_clock),
    .reset(local_pes_9_9_reset),
    .io_in_q(local_pes_9_9_io_in_q),
    .io_in_sum(local_pes_9_9_io_in_sum),
    .io_in_sum_exp(local_pes_9_9_io_in_sum_exp),
    .io_in_kv(local_pes_9_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_9_io_in_inv_sum),
    .io_in_stage(local_pes_9_9_io_in_stage),
    .io_out_q(local_pes_9_9_io_out_q),
    .io_out_sum(local_pes_9_9_io_out_sum),
    .io_out_sum_exp(local_pes_9_9_io_out_sum_exp),
    .io_out_kv(local_pes_9_9_io_out_kv),
    .io_out_stage(local_pes_9_9_io_out_stage)
  );
  PE_1 local_pes_9_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_10_clock),
    .reset(local_pes_9_10_reset),
    .io_in_q(local_pes_9_10_io_in_q),
    .io_in_sum(local_pes_9_10_io_in_sum),
    .io_in_sum_exp(local_pes_9_10_io_in_sum_exp),
    .io_in_kv(local_pes_9_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_10_io_in_inv_sum),
    .io_in_stage(local_pes_9_10_io_in_stage),
    .io_out_q(local_pes_9_10_io_out_q),
    .io_out_sum(local_pes_9_10_io_out_sum),
    .io_out_sum_exp(local_pes_9_10_io_out_sum_exp),
    .io_out_kv(local_pes_9_10_io_out_kv),
    .io_out_stage(local_pes_9_10_io_out_stage)
  );
  PE_1 local_pes_9_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_11_clock),
    .reset(local_pes_9_11_reset),
    .io_in_q(local_pes_9_11_io_in_q),
    .io_in_sum(local_pes_9_11_io_in_sum),
    .io_in_sum_exp(local_pes_9_11_io_in_sum_exp),
    .io_in_kv(local_pes_9_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_11_io_in_inv_sum),
    .io_in_stage(local_pes_9_11_io_in_stage),
    .io_out_q(local_pes_9_11_io_out_q),
    .io_out_sum(local_pes_9_11_io_out_sum),
    .io_out_sum_exp(local_pes_9_11_io_out_sum_exp),
    .io_out_kv(local_pes_9_11_io_out_kv),
    .io_out_stage(local_pes_9_11_io_out_stage)
  );
  PE_1 local_pes_9_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_12_clock),
    .reset(local_pes_9_12_reset),
    .io_in_q(local_pes_9_12_io_in_q),
    .io_in_sum(local_pes_9_12_io_in_sum),
    .io_in_sum_exp(local_pes_9_12_io_in_sum_exp),
    .io_in_kv(local_pes_9_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_12_io_in_inv_sum),
    .io_in_stage(local_pes_9_12_io_in_stage),
    .io_out_q(local_pes_9_12_io_out_q),
    .io_out_sum(local_pes_9_12_io_out_sum),
    .io_out_sum_exp(local_pes_9_12_io_out_sum_exp),
    .io_out_kv(local_pes_9_12_io_out_kv),
    .io_out_stage(local_pes_9_12_io_out_stage)
  );
  PE_1 local_pes_9_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_13_clock),
    .reset(local_pes_9_13_reset),
    .io_in_q(local_pes_9_13_io_in_q),
    .io_in_sum(local_pes_9_13_io_in_sum),
    .io_in_sum_exp(local_pes_9_13_io_in_sum_exp),
    .io_in_kv(local_pes_9_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_13_io_in_inv_sum),
    .io_in_stage(local_pes_9_13_io_in_stage),
    .io_out_q(local_pes_9_13_io_out_q),
    .io_out_sum(local_pes_9_13_io_out_sum),
    .io_out_sum_exp(local_pes_9_13_io_out_sum_exp),
    .io_out_kv(local_pes_9_13_io_out_kv),
    .io_out_stage(local_pes_9_13_io_out_stage)
  );
  PE_1 local_pes_9_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_14_clock),
    .reset(local_pes_9_14_reset),
    .io_in_q(local_pes_9_14_io_in_q),
    .io_in_sum(local_pes_9_14_io_in_sum),
    .io_in_sum_exp(local_pes_9_14_io_in_sum_exp),
    .io_in_kv(local_pes_9_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_14_io_in_inv_sum),
    .io_in_stage(local_pes_9_14_io_in_stage),
    .io_out_q(local_pes_9_14_io_out_q),
    .io_out_sum(local_pes_9_14_io_out_sum),
    .io_out_sum_exp(local_pes_9_14_io_out_sum_exp),
    .io_out_kv(local_pes_9_14_io_out_kv),
    .io_out_stage(local_pes_9_14_io_out_stage)
  );
  PE_1 local_pes_9_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_15_clock),
    .reset(local_pes_9_15_reset),
    .io_in_q(local_pes_9_15_io_in_q),
    .io_in_sum(local_pes_9_15_io_in_sum),
    .io_in_sum_exp(local_pes_9_15_io_in_sum_exp),
    .io_in_kv(local_pes_9_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_15_io_in_inv_sum),
    .io_in_stage(local_pes_9_15_io_in_stage),
    .io_out_q(local_pes_9_15_io_out_q),
    .io_out_sum(local_pes_9_15_io_out_sum),
    .io_out_sum_exp(local_pes_9_15_io_out_sum_exp),
    .io_out_kv(local_pes_9_15_io_out_kv),
    .io_out_stage(local_pes_9_15_io_out_stage)
  );
  PE_1 local_pes_9_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_16_clock),
    .reset(local_pes_9_16_reset),
    .io_in_q(local_pes_9_16_io_in_q),
    .io_in_sum(local_pes_9_16_io_in_sum),
    .io_in_sum_exp(local_pes_9_16_io_in_sum_exp),
    .io_in_kv(local_pes_9_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_16_io_in_inv_sum),
    .io_in_stage(local_pes_9_16_io_in_stage),
    .io_out_q(local_pes_9_16_io_out_q),
    .io_out_sum(local_pes_9_16_io_out_sum),
    .io_out_sum_exp(local_pes_9_16_io_out_sum_exp),
    .io_out_kv(local_pes_9_16_io_out_kv),
    .io_out_stage(local_pes_9_16_io_out_stage)
  );
  PE_1 local_pes_9_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_17_clock),
    .reset(local_pes_9_17_reset),
    .io_in_q(local_pes_9_17_io_in_q),
    .io_in_sum(local_pes_9_17_io_in_sum),
    .io_in_sum_exp(local_pes_9_17_io_in_sum_exp),
    .io_in_kv(local_pes_9_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_17_io_in_inv_sum),
    .io_in_stage(local_pes_9_17_io_in_stage),
    .io_out_q(local_pes_9_17_io_out_q),
    .io_out_sum(local_pes_9_17_io_out_sum),
    .io_out_sum_exp(local_pes_9_17_io_out_sum_exp),
    .io_out_kv(local_pes_9_17_io_out_kv),
    .io_out_stage(local_pes_9_17_io_out_stage)
  );
  PE_1 local_pes_9_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_18_clock),
    .reset(local_pes_9_18_reset),
    .io_in_q(local_pes_9_18_io_in_q),
    .io_in_sum(local_pes_9_18_io_in_sum),
    .io_in_sum_exp(local_pes_9_18_io_in_sum_exp),
    .io_in_kv(local_pes_9_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_18_io_in_inv_sum),
    .io_in_stage(local_pes_9_18_io_in_stage),
    .io_out_q(local_pes_9_18_io_out_q),
    .io_out_sum(local_pes_9_18_io_out_sum),
    .io_out_sum_exp(local_pes_9_18_io_out_sum_exp),
    .io_out_kv(local_pes_9_18_io_out_kv),
    .io_out_stage(local_pes_9_18_io_out_stage)
  );
  PE_1 local_pes_9_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_19_clock),
    .reset(local_pes_9_19_reset),
    .io_in_q(local_pes_9_19_io_in_q),
    .io_in_sum(local_pes_9_19_io_in_sum),
    .io_in_sum_exp(local_pes_9_19_io_in_sum_exp),
    .io_in_kv(local_pes_9_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_19_io_in_inv_sum),
    .io_in_stage(local_pes_9_19_io_in_stage),
    .io_out_q(local_pes_9_19_io_out_q),
    .io_out_sum(local_pes_9_19_io_out_sum),
    .io_out_sum_exp(local_pes_9_19_io_out_sum_exp),
    .io_out_kv(local_pes_9_19_io_out_kv),
    .io_out_stage(local_pes_9_19_io_out_stage)
  );
  PE_1 local_pes_9_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_20_clock),
    .reset(local_pes_9_20_reset),
    .io_in_q(local_pes_9_20_io_in_q),
    .io_in_sum(local_pes_9_20_io_in_sum),
    .io_in_sum_exp(local_pes_9_20_io_in_sum_exp),
    .io_in_kv(local_pes_9_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_20_io_in_inv_sum),
    .io_in_stage(local_pes_9_20_io_in_stage),
    .io_out_q(local_pes_9_20_io_out_q),
    .io_out_sum(local_pes_9_20_io_out_sum),
    .io_out_sum_exp(local_pes_9_20_io_out_sum_exp),
    .io_out_kv(local_pes_9_20_io_out_kv),
    .io_out_stage(local_pes_9_20_io_out_stage)
  );
  PE_1 local_pes_9_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_21_clock),
    .reset(local_pes_9_21_reset),
    .io_in_q(local_pes_9_21_io_in_q),
    .io_in_sum(local_pes_9_21_io_in_sum),
    .io_in_sum_exp(local_pes_9_21_io_in_sum_exp),
    .io_in_kv(local_pes_9_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_21_io_in_inv_sum),
    .io_in_stage(local_pes_9_21_io_in_stage),
    .io_out_q(local_pes_9_21_io_out_q),
    .io_out_sum(local_pes_9_21_io_out_sum),
    .io_out_sum_exp(local_pes_9_21_io_out_sum_exp),
    .io_out_kv(local_pes_9_21_io_out_kv),
    .io_out_stage(local_pes_9_21_io_out_stage)
  );
  PE_1 local_pes_9_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_22_clock),
    .reset(local_pes_9_22_reset),
    .io_in_q(local_pes_9_22_io_in_q),
    .io_in_sum(local_pes_9_22_io_in_sum),
    .io_in_sum_exp(local_pes_9_22_io_in_sum_exp),
    .io_in_kv(local_pes_9_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_22_io_in_inv_sum),
    .io_in_stage(local_pes_9_22_io_in_stage),
    .io_out_q(local_pes_9_22_io_out_q),
    .io_out_sum(local_pes_9_22_io_out_sum),
    .io_out_sum_exp(local_pes_9_22_io_out_sum_exp),
    .io_out_kv(local_pes_9_22_io_out_kv),
    .io_out_stage(local_pes_9_22_io_out_stage)
  );
  PE_1 local_pes_9_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_23_clock),
    .reset(local_pes_9_23_reset),
    .io_in_q(local_pes_9_23_io_in_q),
    .io_in_sum(local_pes_9_23_io_in_sum),
    .io_in_sum_exp(local_pes_9_23_io_in_sum_exp),
    .io_in_kv(local_pes_9_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_23_io_in_inv_sum),
    .io_in_stage(local_pes_9_23_io_in_stage),
    .io_out_q(local_pes_9_23_io_out_q),
    .io_out_sum(local_pes_9_23_io_out_sum),
    .io_out_sum_exp(local_pes_9_23_io_out_sum_exp),
    .io_out_kv(local_pes_9_23_io_out_kv),
    .io_out_stage(local_pes_9_23_io_out_stage)
  );
  PE_1 local_pes_9_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_24_clock),
    .reset(local_pes_9_24_reset),
    .io_in_q(local_pes_9_24_io_in_q),
    .io_in_sum(local_pes_9_24_io_in_sum),
    .io_in_sum_exp(local_pes_9_24_io_in_sum_exp),
    .io_in_kv(local_pes_9_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_24_io_in_inv_sum),
    .io_in_stage(local_pes_9_24_io_in_stage),
    .io_out_q(local_pes_9_24_io_out_q),
    .io_out_sum(local_pes_9_24_io_out_sum),
    .io_out_sum_exp(local_pes_9_24_io_out_sum_exp),
    .io_out_kv(local_pes_9_24_io_out_kv),
    .io_out_stage(local_pes_9_24_io_out_stage)
  );
  PE_1 local_pes_9_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_25_clock),
    .reset(local_pes_9_25_reset),
    .io_in_q(local_pes_9_25_io_in_q),
    .io_in_sum(local_pes_9_25_io_in_sum),
    .io_in_sum_exp(local_pes_9_25_io_in_sum_exp),
    .io_in_kv(local_pes_9_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_25_io_in_inv_sum),
    .io_in_stage(local_pes_9_25_io_in_stage),
    .io_out_q(local_pes_9_25_io_out_q),
    .io_out_sum(local_pes_9_25_io_out_sum),
    .io_out_sum_exp(local_pes_9_25_io_out_sum_exp),
    .io_out_kv(local_pes_9_25_io_out_kv),
    .io_out_stage(local_pes_9_25_io_out_stage)
  );
  PE_1 local_pes_9_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_26_clock),
    .reset(local_pes_9_26_reset),
    .io_in_q(local_pes_9_26_io_in_q),
    .io_in_sum(local_pes_9_26_io_in_sum),
    .io_in_sum_exp(local_pes_9_26_io_in_sum_exp),
    .io_in_kv(local_pes_9_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_26_io_in_inv_sum),
    .io_in_stage(local_pes_9_26_io_in_stage),
    .io_out_q(local_pes_9_26_io_out_q),
    .io_out_sum(local_pes_9_26_io_out_sum),
    .io_out_sum_exp(local_pes_9_26_io_out_sum_exp),
    .io_out_kv(local_pes_9_26_io_out_kv),
    .io_out_stage(local_pes_9_26_io_out_stage)
  );
  PE_1 local_pes_9_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_27_clock),
    .reset(local_pes_9_27_reset),
    .io_in_q(local_pes_9_27_io_in_q),
    .io_in_sum(local_pes_9_27_io_in_sum),
    .io_in_sum_exp(local_pes_9_27_io_in_sum_exp),
    .io_in_kv(local_pes_9_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_27_io_in_inv_sum),
    .io_in_stage(local_pes_9_27_io_in_stage),
    .io_out_q(local_pes_9_27_io_out_q),
    .io_out_sum(local_pes_9_27_io_out_sum),
    .io_out_sum_exp(local_pes_9_27_io_out_sum_exp),
    .io_out_kv(local_pes_9_27_io_out_kv),
    .io_out_stage(local_pes_9_27_io_out_stage)
  );
  PE_1 local_pes_9_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_28_clock),
    .reset(local_pes_9_28_reset),
    .io_in_q(local_pes_9_28_io_in_q),
    .io_in_sum(local_pes_9_28_io_in_sum),
    .io_in_sum_exp(local_pes_9_28_io_in_sum_exp),
    .io_in_kv(local_pes_9_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_28_io_in_inv_sum),
    .io_in_stage(local_pes_9_28_io_in_stage),
    .io_out_q(local_pes_9_28_io_out_q),
    .io_out_sum(local_pes_9_28_io_out_sum),
    .io_out_sum_exp(local_pes_9_28_io_out_sum_exp),
    .io_out_kv(local_pes_9_28_io_out_kv),
    .io_out_stage(local_pes_9_28_io_out_stage)
  );
  PE_1 local_pes_9_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_29_clock),
    .reset(local_pes_9_29_reset),
    .io_in_q(local_pes_9_29_io_in_q),
    .io_in_sum(local_pes_9_29_io_in_sum),
    .io_in_sum_exp(local_pes_9_29_io_in_sum_exp),
    .io_in_kv(local_pes_9_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_29_io_in_inv_sum),
    .io_in_stage(local_pes_9_29_io_in_stage),
    .io_out_q(local_pes_9_29_io_out_q),
    .io_out_sum(local_pes_9_29_io_out_sum),
    .io_out_sum_exp(local_pes_9_29_io_out_sum_exp),
    .io_out_kv(local_pes_9_29_io_out_kv),
    .io_out_stage(local_pes_9_29_io_out_stage)
  );
  PE_1 local_pes_9_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_30_clock),
    .reset(local_pes_9_30_reset),
    .io_in_q(local_pes_9_30_io_in_q),
    .io_in_sum(local_pes_9_30_io_in_sum),
    .io_in_sum_exp(local_pes_9_30_io_in_sum_exp),
    .io_in_kv(local_pes_9_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_30_io_in_inv_sum),
    .io_in_stage(local_pes_9_30_io_in_stage),
    .io_out_q(local_pes_9_30_io_out_q),
    .io_out_sum(local_pes_9_30_io_out_sum),
    .io_out_sum_exp(local_pes_9_30_io_out_sum_exp),
    .io_out_kv(local_pes_9_30_io_out_kv),
    .io_out_stage(local_pes_9_30_io_out_stage)
  );
  PE_1 local_pes_9_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_9_31_clock),
    .reset(local_pes_9_31_reset),
    .io_in_q(local_pes_9_31_io_in_q),
    .io_in_sum(local_pes_9_31_io_in_sum),
    .io_in_sum_exp(local_pes_9_31_io_in_sum_exp),
    .io_in_kv(local_pes_9_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_9_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_9_31_io_in_inv_sum),
    .io_in_stage(local_pes_9_31_io_in_stage),
    .io_out_q(local_pes_9_31_io_out_q),
    .io_out_sum(local_pes_9_31_io_out_sum),
    .io_out_sum_exp(local_pes_9_31_io_out_sum_exp),
    .io_out_kv(local_pes_9_31_io_out_kv),
    .io_out_stage(local_pes_9_31_io_out_stage)
  );
  PE local_pes_10_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_0_clock),
    .reset(local_pes_10_0_reset),
    .io_in_q(local_pes_10_0_io_in_q),
    .io_in_kv(local_pes_10_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_0_io_in_inv_sum),
    .io_in_stage(local_pes_10_0_io_in_stage),
    .io_out_q(local_pes_10_0_io_out_q),
    .io_out_sum(local_pes_10_0_io_out_sum),
    .io_out_kv(local_pes_10_0_io_out_kv),
    .io_out_stage(local_pes_10_0_io_out_stage)
  );
  PE_1 local_pes_10_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_1_clock),
    .reset(local_pes_10_1_reset),
    .io_in_q(local_pes_10_1_io_in_q),
    .io_in_sum(local_pes_10_1_io_in_sum),
    .io_in_sum_exp(local_pes_10_1_io_in_sum_exp),
    .io_in_kv(local_pes_10_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_1_io_in_inv_sum),
    .io_in_stage(local_pes_10_1_io_in_stage),
    .io_out_q(local_pes_10_1_io_out_q),
    .io_out_sum(local_pes_10_1_io_out_sum),
    .io_out_sum_exp(local_pes_10_1_io_out_sum_exp),
    .io_out_kv(local_pes_10_1_io_out_kv),
    .io_out_stage(local_pes_10_1_io_out_stage)
  );
  PE_1 local_pes_10_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_2_clock),
    .reset(local_pes_10_2_reset),
    .io_in_q(local_pes_10_2_io_in_q),
    .io_in_sum(local_pes_10_2_io_in_sum),
    .io_in_sum_exp(local_pes_10_2_io_in_sum_exp),
    .io_in_kv(local_pes_10_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_2_io_in_inv_sum),
    .io_in_stage(local_pes_10_2_io_in_stage),
    .io_out_q(local_pes_10_2_io_out_q),
    .io_out_sum(local_pes_10_2_io_out_sum),
    .io_out_sum_exp(local_pes_10_2_io_out_sum_exp),
    .io_out_kv(local_pes_10_2_io_out_kv),
    .io_out_stage(local_pes_10_2_io_out_stage)
  );
  PE_1 local_pes_10_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_3_clock),
    .reset(local_pes_10_3_reset),
    .io_in_q(local_pes_10_3_io_in_q),
    .io_in_sum(local_pes_10_3_io_in_sum),
    .io_in_sum_exp(local_pes_10_3_io_in_sum_exp),
    .io_in_kv(local_pes_10_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_3_io_in_inv_sum),
    .io_in_stage(local_pes_10_3_io_in_stage),
    .io_out_q(local_pes_10_3_io_out_q),
    .io_out_sum(local_pes_10_3_io_out_sum),
    .io_out_sum_exp(local_pes_10_3_io_out_sum_exp),
    .io_out_kv(local_pes_10_3_io_out_kv),
    .io_out_stage(local_pes_10_3_io_out_stage)
  );
  PE_1 local_pes_10_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_4_clock),
    .reset(local_pes_10_4_reset),
    .io_in_q(local_pes_10_4_io_in_q),
    .io_in_sum(local_pes_10_4_io_in_sum),
    .io_in_sum_exp(local_pes_10_4_io_in_sum_exp),
    .io_in_kv(local_pes_10_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_4_io_in_inv_sum),
    .io_in_stage(local_pes_10_4_io_in_stage),
    .io_out_q(local_pes_10_4_io_out_q),
    .io_out_sum(local_pes_10_4_io_out_sum),
    .io_out_sum_exp(local_pes_10_4_io_out_sum_exp),
    .io_out_kv(local_pes_10_4_io_out_kv),
    .io_out_stage(local_pes_10_4_io_out_stage)
  );
  PE_1 local_pes_10_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_5_clock),
    .reset(local_pes_10_5_reset),
    .io_in_q(local_pes_10_5_io_in_q),
    .io_in_sum(local_pes_10_5_io_in_sum),
    .io_in_sum_exp(local_pes_10_5_io_in_sum_exp),
    .io_in_kv(local_pes_10_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_5_io_in_inv_sum),
    .io_in_stage(local_pes_10_5_io_in_stage),
    .io_out_q(local_pes_10_5_io_out_q),
    .io_out_sum(local_pes_10_5_io_out_sum),
    .io_out_sum_exp(local_pes_10_5_io_out_sum_exp),
    .io_out_kv(local_pes_10_5_io_out_kv),
    .io_out_stage(local_pes_10_5_io_out_stage)
  );
  PE_1 local_pes_10_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_6_clock),
    .reset(local_pes_10_6_reset),
    .io_in_q(local_pes_10_6_io_in_q),
    .io_in_sum(local_pes_10_6_io_in_sum),
    .io_in_sum_exp(local_pes_10_6_io_in_sum_exp),
    .io_in_kv(local_pes_10_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_6_io_in_inv_sum),
    .io_in_stage(local_pes_10_6_io_in_stage),
    .io_out_q(local_pes_10_6_io_out_q),
    .io_out_sum(local_pes_10_6_io_out_sum),
    .io_out_sum_exp(local_pes_10_6_io_out_sum_exp),
    .io_out_kv(local_pes_10_6_io_out_kv),
    .io_out_stage(local_pes_10_6_io_out_stage)
  );
  PE_1 local_pes_10_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_7_clock),
    .reset(local_pes_10_7_reset),
    .io_in_q(local_pes_10_7_io_in_q),
    .io_in_sum(local_pes_10_7_io_in_sum),
    .io_in_sum_exp(local_pes_10_7_io_in_sum_exp),
    .io_in_kv(local_pes_10_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_7_io_in_inv_sum),
    .io_in_stage(local_pes_10_7_io_in_stage),
    .io_out_q(local_pes_10_7_io_out_q),
    .io_out_sum(local_pes_10_7_io_out_sum),
    .io_out_sum_exp(local_pes_10_7_io_out_sum_exp),
    .io_out_kv(local_pes_10_7_io_out_kv),
    .io_out_stage(local_pes_10_7_io_out_stage)
  );
  PE_1 local_pes_10_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_8_clock),
    .reset(local_pes_10_8_reset),
    .io_in_q(local_pes_10_8_io_in_q),
    .io_in_sum(local_pes_10_8_io_in_sum),
    .io_in_sum_exp(local_pes_10_8_io_in_sum_exp),
    .io_in_kv(local_pes_10_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_8_io_in_inv_sum),
    .io_in_stage(local_pes_10_8_io_in_stage),
    .io_out_q(local_pes_10_8_io_out_q),
    .io_out_sum(local_pes_10_8_io_out_sum),
    .io_out_sum_exp(local_pes_10_8_io_out_sum_exp),
    .io_out_kv(local_pes_10_8_io_out_kv),
    .io_out_stage(local_pes_10_8_io_out_stage)
  );
  PE_1 local_pes_10_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_9_clock),
    .reset(local_pes_10_9_reset),
    .io_in_q(local_pes_10_9_io_in_q),
    .io_in_sum(local_pes_10_9_io_in_sum),
    .io_in_sum_exp(local_pes_10_9_io_in_sum_exp),
    .io_in_kv(local_pes_10_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_9_io_in_inv_sum),
    .io_in_stage(local_pes_10_9_io_in_stage),
    .io_out_q(local_pes_10_9_io_out_q),
    .io_out_sum(local_pes_10_9_io_out_sum),
    .io_out_sum_exp(local_pes_10_9_io_out_sum_exp),
    .io_out_kv(local_pes_10_9_io_out_kv),
    .io_out_stage(local_pes_10_9_io_out_stage)
  );
  PE_1 local_pes_10_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_10_clock),
    .reset(local_pes_10_10_reset),
    .io_in_q(local_pes_10_10_io_in_q),
    .io_in_sum(local_pes_10_10_io_in_sum),
    .io_in_sum_exp(local_pes_10_10_io_in_sum_exp),
    .io_in_kv(local_pes_10_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_10_io_in_inv_sum),
    .io_in_stage(local_pes_10_10_io_in_stage),
    .io_out_q(local_pes_10_10_io_out_q),
    .io_out_sum(local_pes_10_10_io_out_sum),
    .io_out_sum_exp(local_pes_10_10_io_out_sum_exp),
    .io_out_kv(local_pes_10_10_io_out_kv),
    .io_out_stage(local_pes_10_10_io_out_stage)
  );
  PE_1 local_pes_10_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_11_clock),
    .reset(local_pes_10_11_reset),
    .io_in_q(local_pes_10_11_io_in_q),
    .io_in_sum(local_pes_10_11_io_in_sum),
    .io_in_sum_exp(local_pes_10_11_io_in_sum_exp),
    .io_in_kv(local_pes_10_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_11_io_in_inv_sum),
    .io_in_stage(local_pes_10_11_io_in_stage),
    .io_out_q(local_pes_10_11_io_out_q),
    .io_out_sum(local_pes_10_11_io_out_sum),
    .io_out_sum_exp(local_pes_10_11_io_out_sum_exp),
    .io_out_kv(local_pes_10_11_io_out_kv),
    .io_out_stage(local_pes_10_11_io_out_stage)
  );
  PE_1 local_pes_10_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_12_clock),
    .reset(local_pes_10_12_reset),
    .io_in_q(local_pes_10_12_io_in_q),
    .io_in_sum(local_pes_10_12_io_in_sum),
    .io_in_sum_exp(local_pes_10_12_io_in_sum_exp),
    .io_in_kv(local_pes_10_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_12_io_in_inv_sum),
    .io_in_stage(local_pes_10_12_io_in_stage),
    .io_out_q(local_pes_10_12_io_out_q),
    .io_out_sum(local_pes_10_12_io_out_sum),
    .io_out_sum_exp(local_pes_10_12_io_out_sum_exp),
    .io_out_kv(local_pes_10_12_io_out_kv),
    .io_out_stage(local_pes_10_12_io_out_stage)
  );
  PE_1 local_pes_10_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_13_clock),
    .reset(local_pes_10_13_reset),
    .io_in_q(local_pes_10_13_io_in_q),
    .io_in_sum(local_pes_10_13_io_in_sum),
    .io_in_sum_exp(local_pes_10_13_io_in_sum_exp),
    .io_in_kv(local_pes_10_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_13_io_in_inv_sum),
    .io_in_stage(local_pes_10_13_io_in_stage),
    .io_out_q(local_pes_10_13_io_out_q),
    .io_out_sum(local_pes_10_13_io_out_sum),
    .io_out_sum_exp(local_pes_10_13_io_out_sum_exp),
    .io_out_kv(local_pes_10_13_io_out_kv),
    .io_out_stage(local_pes_10_13_io_out_stage)
  );
  PE_1 local_pes_10_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_14_clock),
    .reset(local_pes_10_14_reset),
    .io_in_q(local_pes_10_14_io_in_q),
    .io_in_sum(local_pes_10_14_io_in_sum),
    .io_in_sum_exp(local_pes_10_14_io_in_sum_exp),
    .io_in_kv(local_pes_10_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_14_io_in_inv_sum),
    .io_in_stage(local_pes_10_14_io_in_stage),
    .io_out_q(local_pes_10_14_io_out_q),
    .io_out_sum(local_pes_10_14_io_out_sum),
    .io_out_sum_exp(local_pes_10_14_io_out_sum_exp),
    .io_out_kv(local_pes_10_14_io_out_kv),
    .io_out_stage(local_pes_10_14_io_out_stage)
  );
  PE_1 local_pes_10_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_15_clock),
    .reset(local_pes_10_15_reset),
    .io_in_q(local_pes_10_15_io_in_q),
    .io_in_sum(local_pes_10_15_io_in_sum),
    .io_in_sum_exp(local_pes_10_15_io_in_sum_exp),
    .io_in_kv(local_pes_10_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_15_io_in_inv_sum),
    .io_in_stage(local_pes_10_15_io_in_stage),
    .io_out_q(local_pes_10_15_io_out_q),
    .io_out_sum(local_pes_10_15_io_out_sum),
    .io_out_sum_exp(local_pes_10_15_io_out_sum_exp),
    .io_out_kv(local_pes_10_15_io_out_kv),
    .io_out_stage(local_pes_10_15_io_out_stage)
  );
  PE_1 local_pes_10_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_16_clock),
    .reset(local_pes_10_16_reset),
    .io_in_q(local_pes_10_16_io_in_q),
    .io_in_sum(local_pes_10_16_io_in_sum),
    .io_in_sum_exp(local_pes_10_16_io_in_sum_exp),
    .io_in_kv(local_pes_10_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_16_io_in_inv_sum),
    .io_in_stage(local_pes_10_16_io_in_stage),
    .io_out_q(local_pes_10_16_io_out_q),
    .io_out_sum(local_pes_10_16_io_out_sum),
    .io_out_sum_exp(local_pes_10_16_io_out_sum_exp),
    .io_out_kv(local_pes_10_16_io_out_kv),
    .io_out_stage(local_pes_10_16_io_out_stage)
  );
  PE_1 local_pes_10_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_17_clock),
    .reset(local_pes_10_17_reset),
    .io_in_q(local_pes_10_17_io_in_q),
    .io_in_sum(local_pes_10_17_io_in_sum),
    .io_in_sum_exp(local_pes_10_17_io_in_sum_exp),
    .io_in_kv(local_pes_10_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_17_io_in_inv_sum),
    .io_in_stage(local_pes_10_17_io_in_stage),
    .io_out_q(local_pes_10_17_io_out_q),
    .io_out_sum(local_pes_10_17_io_out_sum),
    .io_out_sum_exp(local_pes_10_17_io_out_sum_exp),
    .io_out_kv(local_pes_10_17_io_out_kv),
    .io_out_stage(local_pes_10_17_io_out_stage)
  );
  PE_1 local_pes_10_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_18_clock),
    .reset(local_pes_10_18_reset),
    .io_in_q(local_pes_10_18_io_in_q),
    .io_in_sum(local_pes_10_18_io_in_sum),
    .io_in_sum_exp(local_pes_10_18_io_in_sum_exp),
    .io_in_kv(local_pes_10_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_18_io_in_inv_sum),
    .io_in_stage(local_pes_10_18_io_in_stage),
    .io_out_q(local_pes_10_18_io_out_q),
    .io_out_sum(local_pes_10_18_io_out_sum),
    .io_out_sum_exp(local_pes_10_18_io_out_sum_exp),
    .io_out_kv(local_pes_10_18_io_out_kv),
    .io_out_stage(local_pes_10_18_io_out_stage)
  );
  PE_1 local_pes_10_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_19_clock),
    .reset(local_pes_10_19_reset),
    .io_in_q(local_pes_10_19_io_in_q),
    .io_in_sum(local_pes_10_19_io_in_sum),
    .io_in_sum_exp(local_pes_10_19_io_in_sum_exp),
    .io_in_kv(local_pes_10_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_19_io_in_inv_sum),
    .io_in_stage(local_pes_10_19_io_in_stage),
    .io_out_q(local_pes_10_19_io_out_q),
    .io_out_sum(local_pes_10_19_io_out_sum),
    .io_out_sum_exp(local_pes_10_19_io_out_sum_exp),
    .io_out_kv(local_pes_10_19_io_out_kv),
    .io_out_stage(local_pes_10_19_io_out_stage)
  );
  PE_1 local_pes_10_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_20_clock),
    .reset(local_pes_10_20_reset),
    .io_in_q(local_pes_10_20_io_in_q),
    .io_in_sum(local_pes_10_20_io_in_sum),
    .io_in_sum_exp(local_pes_10_20_io_in_sum_exp),
    .io_in_kv(local_pes_10_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_20_io_in_inv_sum),
    .io_in_stage(local_pes_10_20_io_in_stage),
    .io_out_q(local_pes_10_20_io_out_q),
    .io_out_sum(local_pes_10_20_io_out_sum),
    .io_out_sum_exp(local_pes_10_20_io_out_sum_exp),
    .io_out_kv(local_pes_10_20_io_out_kv),
    .io_out_stage(local_pes_10_20_io_out_stage)
  );
  PE_1 local_pes_10_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_21_clock),
    .reset(local_pes_10_21_reset),
    .io_in_q(local_pes_10_21_io_in_q),
    .io_in_sum(local_pes_10_21_io_in_sum),
    .io_in_sum_exp(local_pes_10_21_io_in_sum_exp),
    .io_in_kv(local_pes_10_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_21_io_in_inv_sum),
    .io_in_stage(local_pes_10_21_io_in_stage),
    .io_out_q(local_pes_10_21_io_out_q),
    .io_out_sum(local_pes_10_21_io_out_sum),
    .io_out_sum_exp(local_pes_10_21_io_out_sum_exp),
    .io_out_kv(local_pes_10_21_io_out_kv),
    .io_out_stage(local_pes_10_21_io_out_stage)
  );
  PE_1 local_pes_10_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_22_clock),
    .reset(local_pes_10_22_reset),
    .io_in_q(local_pes_10_22_io_in_q),
    .io_in_sum(local_pes_10_22_io_in_sum),
    .io_in_sum_exp(local_pes_10_22_io_in_sum_exp),
    .io_in_kv(local_pes_10_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_22_io_in_inv_sum),
    .io_in_stage(local_pes_10_22_io_in_stage),
    .io_out_q(local_pes_10_22_io_out_q),
    .io_out_sum(local_pes_10_22_io_out_sum),
    .io_out_sum_exp(local_pes_10_22_io_out_sum_exp),
    .io_out_kv(local_pes_10_22_io_out_kv),
    .io_out_stage(local_pes_10_22_io_out_stage)
  );
  PE_1 local_pes_10_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_23_clock),
    .reset(local_pes_10_23_reset),
    .io_in_q(local_pes_10_23_io_in_q),
    .io_in_sum(local_pes_10_23_io_in_sum),
    .io_in_sum_exp(local_pes_10_23_io_in_sum_exp),
    .io_in_kv(local_pes_10_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_23_io_in_inv_sum),
    .io_in_stage(local_pes_10_23_io_in_stage),
    .io_out_q(local_pes_10_23_io_out_q),
    .io_out_sum(local_pes_10_23_io_out_sum),
    .io_out_sum_exp(local_pes_10_23_io_out_sum_exp),
    .io_out_kv(local_pes_10_23_io_out_kv),
    .io_out_stage(local_pes_10_23_io_out_stage)
  );
  PE_1 local_pes_10_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_24_clock),
    .reset(local_pes_10_24_reset),
    .io_in_q(local_pes_10_24_io_in_q),
    .io_in_sum(local_pes_10_24_io_in_sum),
    .io_in_sum_exp(local_pes_10_24_io_in_sum_exp),
    .io_in_kv(local_pes_10_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_24_io_in_inv_sum),
    .io_in_stage(local_pes_10_24_io_in_stage),
    .io_out_q(local_pes_10_24_io_out_q),
    .io_out_sum(local_pes_10_24_io_out_sum),
    .io_out_sum_exp(local_pes_10_24_io_out_sum_exp),
    .io_out_kv(local_pes_10_24_io_out_kv),
    .io_out_stage(local_pes_10_24_io_out_stage)
  );
  PE_1 local_pes_10_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_25_clock),
    .reset(local_pes_10_25_reset),
    .io_in_q(local_pes_10_25_io_in_q),
    .io_in_sum(local_pes_10_25_io_in_sum),
    .io_in_sum_exp(local_pes_10_25_io_in_sum_exp),
    .io_in_kv(local_pes_10_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_25_io_in_inv_sum),
    .io_in_stage(local_pes_10_25_io_in_stage),
    .io_out_q(local_pes_10_25_io_out_q),
    .io_out_sum(local_pes_10_25_io_out_sum),
    .io_out_sum_exp(local_pes_10_25_io_out_sum_exp),
    .io_out_kv(local_pes_10_25_io_out_kv),
    .io_out_stage(local_pes_10_25_io_out_stage)
  );
  PE_1 local_pes_10_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_26_clock),
    .reset(local_pes_10_26_reset),
    .io_in_q(local_pes_10_26_io_in_q),
    .io_in_sum(local_pes_10_26_io_in_sum),
    .io_in_sum_exp(local_pes_10_26_io_in_sum_exp),
    .io_in_kv(local_pes_10_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_26_io_in_inv_sum),
    .io_in_stage(local_pes_10_26_io_in_stage),
    .io_out_q(local_pes_10_26_io_out_q),
    .io_out_sum(local_pes_10_26_io_out_sum),
    .io_out_sum_exp(local_pes_10_26_io_out_sum_exp),
    .io_out_kv(local_pes_10_26_io_out_kv),
    .io_out_stage(local_pes_10_26_io_out_stage)
  );
  PE_1 local_pes_10_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_27_clock),
    .reset(local_pes_10_27_reset),
    .io_in_q(local_pes_10_27_io_in_q),
    .io_in_sum(local_pes_10_27_io_in_sum),
    .io_in_sum_exp(local_pes_10_27_io_in_sum_exp),
    .io_in_kv(local_pes_10_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_27_io_in_inv_sum),
    .io_in_stage(local_pes_10_27_io_in_stage),
    .io_out_q(local_pes_10_27_io_out_q),
    .io_out_sum(local_pes_10_27_io_out_sum),
    .io_out_sum_exp(local_pes_10_27_io_out_sum_exp),
    .io_out_kv(local_pes_10_27_io_out_kv),
    .io_out_stage(local_pes_10_27_io_out_stage)
  );
  PE_1 local_pes_10_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_28_clock),
    .reset(local_pes_10_28_reset),
    .io_in_q(local_pes_10_28_io_in_q),
    .io_in_sum(local_pes_10_28_io_in_sum),
    .io_in_sum_exp(local_pes_10_28_io_in_sum_exp),
    .io_in_kv(local_pes_10_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_28_io_in_inv_sum),
    .io_in_stage(local_pes_10_28_io_in_stage),
    .io_out_q(local_pes_10_28_io_out_q),
    .io_out_sum(local_pes_10_28_io_out_sum),
    .io_out_sum_exp(local_pes_10_28_io_out_sum_exp),
    .io_out_kv(local_pes_10_28_io_out_kv),
    .io_out_stage(local_pes_10_28_io_out_stage)
  );
  PE_1 local_pes_10_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_29_clock),
    .reset(local_pes_10_29_reset),
    .io_in_q(local_pes_10_29_io_in_q),
    .io_in_sum(local_pes_10_29_io_in_sum),
    .io_in_sum_exp(local_pes_10_29_io_in_sum_exp),
    .io_in_kv(local_pes_10_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_29_io_in_inv_sum),
    .io_in_stage(local_pes_10_29_io_in_stage),
    .io_out_q(local_pes_10_29_io_out_q),
    .io_out_sum(local_pes_10_29_io_out_sum),
    .io_out_sum_exp(local_pes_10_29_io_out_sum_exp),
    .io_out_kv(local_pes_10_29_io_out_kv),
    .io_out_stage(local_pes_10_29_io_out_stage)
  );
  PE_1 local_pes_10_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_30_clock),
    .reset(local_pes_10_30_reset),
    .io_in_q(local_pes_10_30_io_in_q),
    .io_in_sum(local_pes_10_30_io_in_sum),
    .io_in_sum_exp(local_pes_10_30_io_in_sum_exp),
    .io_in_kv(local_pes_10_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_30_io_in_inv_sum),
    .io_in_stage(local_pes_10_30_io_in_stage),
    .io_out_q(local_pes_10_30_io_out_q),
    .io_out_sum(local_pes_10_30_io_out_sum),
    .io_out_sum_exp(local_pes_10_30_io_out_sum_exp),
    .io_out_kv(local_pes_10_30_io_out_kv),
    .io_out_stage(local_pes_10_30_io_out_stage)
  );
  PE_1 local_pes_10_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_10_31_clock),
    .reset(local_pes_10_31_reset),
    .io_in_q(local_pes_10_31_io_in_q),
    .io_in_sum(local_pes_10_31_io_in_sum),
    .io_in_sum_exp(local_pes_10_31_io_in_sum_exp),
    .io_in_kv(local_pes_10_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_10_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_10_31_io_in_inv_sum),
    .io_in_stage(local_pes_10_31_io_in_stage),
    .io_out_q(local_pes_10_31_io_out_q),
    .io_out_sum(local_pes_10_31_io_out_sum),
    .io_out_sum_exp(local_pes_10_31_io_out_sum_exp),
    .io_out_kv(local_pes_10_31_io_out_kv),
    .io_out_stage(local_pes_10_31_io_out_stage)
  );
  PE local_pes_11_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_0_clock),
    .reset(local_pes_11_0_reset),
    .io_in_q(local_pes_11_0_io_in_q),
    .io_in_kv(local_pes_11_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_0_io_in_inv_sum),
    .io_in_stage(local_pes_11_0_io_in_stage),
    .io_out_q(local_pes_11_0_io_out_q),
    .io_out_sum(local_pes_11_0_io_out_sum),
    .io_out_kv(local_pes_11_0_io_out_kv),
    .io_out_stage(local_pes_11_0_io_out_stage)
  );
  PE_1 local_pes_11_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_1_clock),
    .reset(local_pes_11_1_reset),
    .io_in_q(local_pes_11_1_io_in_q),
    .io_in_sum(local_pes_11_1_io_in_sum),
    .io_in_sum_exp(local_pes_11_1_io_in_sum_exp),
    .io_in_kv(local_pes_11_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_1_io_in_inv_sum),
    .io_in_stage(local_pes_11_1_io_in_stage),
    .io_out_q(local_pes_11_1_io_out_q),
    .io_out_sum(local_pes_11_1_io_out_sum),
    .io_out_sum_exp(local_pes_11_1_io_out_sum_exp),
    .io_out_kv(local_pes_11_1_io_out_kv),
    .io_out_stage(local_pes_11_1_io_out_stage)
  );
  PE_1 local_pes_11_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_2_clock),
    .reset(local_pes_11_2_reset),
    .io_in_q(local_pes_11_2_io_in_q),
    .io_in_sum(local_pes_11_2_io_in_sum),
    .io_in_sum_exp(local_pes_11_2_io_in_sum_exp),
    .io_in_kv(local_pes_11_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_2_io_in_inv_sum),
    .io_in_stage(local_pes_11_2_io_in_stage),
    .io_out_q(local_pes_11_2_io_out_q),
    .io_out_sum(local_pes_11_2_io_out_sum),
    .io_out_sum_exp(local_pes_11_2_io_out_sum_exp),
    .io_out_kv(local_pes_11_2_io_out_kv),
    .io_out_stage(local_pes_11_2_io_out_stage)
  );
  PE_1 local_pes_11_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_3_clock),
    .reset(local_pes_11_3_reset),
    .io_in_q(local_pes_11_3_io_in_q),
    .io_in_sum(local_pes_11_3_io_in_sum),
    .io_in_sum_exp(local_pes_11_3_io_in_sum_exp),
    .io_in_kv(local_pes_11_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_3_io_in_inv_sum),
    .io_in_stage(local_pes_11_3_io_in_stage),
    .io_out_q(local_pes_11_3_io_out_q),
    .io_out_sum(local_pes_11_3_io_out_sum),
    .io_out_sum_exp(local_pes_11_3_io_out_sum_exp),
    .io_out_kv(local_pes_11_3_io_out_kv),
    .io_out_stage(local_pes_11_3_io_out_stage)
  );
  PE_1 local_pes_11_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_4_clock),
    .reset(local_pes_11_4_reset),
    .io_in_q(local_pes_11_4_io_in_q),
    .io_in_sum(local_pes_11_4_io_in_sum),
    .io_in_sum_exp(local_pes_11_4_io_in_sum_exp),
    .io_in_kv(local_pes_11_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_4_io_in_inv_sum),
    .io_in_stage(local_pes_11_4_io_in_stage),
    .io_out_q(local_pes_11_4_io_out_q),
    .io_out_sum(local_pes_11_4_io_out_sum),
    .io_out_sum_exp(local_pes_11_4_io_out_sum_exp),
    .io_out_kv(local_pes_11_4_io_out_kv),
    .io_out_stage(local_pes_11_4_io_out_stage)
  );
  PE_1 local_pes_11_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_5_clock),
    .reset(local_pes_11_5_reset),
    .io_in_q(local_pes_11_5_io_in_q),
    .io_in_sum(local_pes_11_5_io_in_sum),
    .io_in_sum_exp(local_pes_11_5_io_in_sum_exp),
    .io_in_kv(local_pes_11_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_5_io_in_inv_sum),
    .io_in_stage(local_pes_11_5_io_in_stage),
    .io_out_q(local_pes_11_5_io_out_q),
    .io_out_sum(local_pes_11_5_io_out_sum),
    .io_out_sum_exp(local_pes_11_5_io_out_sum_exp),
    .io_out_kv(local_pes_11_5_io_out_kv),
    .io_out_stage(local_pes_11_5_io_out_stage)
  );
  PE_1 local_pes_11_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_6_clock),
    .reset(local_pes_11_6_reset),
    .io_in_q(local_pes_11_6_io_in_q),
    .io_in_sum(local_pes_11_6_io_in_sum),
    .io_in_sum_exp(local_pes_11_6_io_in_sum_exp),
    .io_in_kv(local_pes_11_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_6_io_in_inv_sum),
    .io_in_stage(local_pes_11_6_io_in_stage),
    .io_out_q(local_pes_11_6_io_out_q),
    .io_out_sum(local_pes_11_6_io_out_sum),
    .io_out_sum_exp(local_pes_11_6_io_out_sum_exp),
    .io_out_kv(local_pes_11_6_io_out_kv),
    .io_out_stage(local_pes_11_6_io_out_stage)
  );
  PE_1 local_pes_11_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_7_clock),
    .reset(local_pes_11_7_reset),
    .io_in_q(local_pes_11_7_io_in_q),
    .io_in_sum(local_pes_11_7_io_in_sum),
    .io_in_sum_exp(local_pes_11_7_io_in_sum_exp),
    .io_in_kv(local_pes_11_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_7_io_in_inv_sum),
    .io_in_stage(local_pes_11_7_io_in_stage),
    .io_out_q(local_pes_11_7_io_out_q),
    .io_out_sum(local_pes_11_7_io_out_sum),
    .io_out_sum_exp(local_pes_11_7_io_out_sum_exp),
    .io_out_kv(local_pes_11_7_io_out_kv),
    .io_out_stage(local_pes_11_7_io_out_stage)
  );
  PE_1 local_pes_11_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_8_clock),
    .reset(local_pes_11_8_reset),
    .io_in_q(local_pes_11_8_io_in_q),
    .io_in_sum(local_pes_11_8_io_in_sum),
    .io_in_sum_exp(local_pes_11_8_io_in_sum_exp),
    .io_in_kv(local_pes_11_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_8_io_in_inv_sum),
    .io_in_stage(local_pes_11_8_io_in_stage),
    .io_out_q(local_pes_11_8_io_out_q),
    .io_out_sum(local_pes_11_8_io_out_sum),
    .io_out_sum_exp(local_pes_11_8_io_out_sum_exp),
    .io_out_kv(local_pes_11_8_io_out_kv),
    .io_out_stage(local_pes_11_8_io_out_stage)
  );
  PE_1 local_pes_11_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_9_clock),
    .reset(local_pes_11_9_reset),
    .io_in_q(local_pes_11_9_io_in_q),
    .io_in_sum(local_pes_11_9_io_in_sum),
    .io_in_sum_exp(local_pes_11_9_io_in_sum_exp),
    .io_in_kv(local_pes_11_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_9_io_in_inv_sum),
    .io_in_stage(local_pes_11_9_io_in_stage),
    .io_out_q(local_pes_11_9_io_out_q),
    .io_out_sum(local_pes_11_9_io_out_sum),
    .io_out_sum_exp(local_pes_11_9_io_out_sum_exp),
    .io_out_kv(local_pes_11_9_io_out_kv),
    .io_out_stage(local_pes_11_9_io_out_stage)
  );
  PE_1 local_pes_11_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_10_clock),
    .reset(local_pes_11_10_reset),
    .io_in_q(local_pes_11_10_io_in_q),
    .io_in_sum(local_pes_11_10_io_in_sum),
    .io_in_sum_exp(local_pes_11_10_io_in_sum_exp),
    .io_in_kv(local_pes_11_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_10_io_in_inv_sum),
    .io_in_stage(local_pes_11_10_io_in_stage),
    .io_out_q(local_pes_11_10_io_out_q),
    .io_out_sum(local_pes_11_10_io_out_sum),
    .io_out_sum_exp(local_pes_11_10_io_out_sum_exp),
    .io_out_kv(local_pes_11_10_io_out_kv),
    .io_out_stage(local_pes_11_10_io_out_stage)
  );
  PE_1 local_pes_11_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_11_clock),
    .reset(local_pes_11_11_reset),
    .io_in_q(local_pes_11_11_io_in_q),
    .io_in_sum(local_pes_11_11_io_in_sum),
    .io_in_sum_exp(local_pes_11_11_io_in_sum_exp),
    .io_in_kv(local_pes_11_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_11_io_in_inv_sum),
    .io_in_stage(local_pes_11_11_io_in_stage),
    .io_out_q(local_pes_11_11_io_out_q),
    .io_out_sum(local_pes_11_11_io_out_sum),
    .io_out_sum_exp(local_pes_11_11_io_out_sum_exp),
    .io_out_kv(local_pes_11_11_io_out_kv),
    .io_out_stage(local_pes_11_11_io_out_stage)
  );
  PE_1 local_pes_11_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_12_clock),
    .reset(local_pes_11_12_reset),
    .io_in_q(local_pes_11_12_io_in_q),
    .io_in_sum(local_pes_11_12_io_in_sum),
    .io_in_sum_exp(local_pes_11_12_io_in_sum_exp),
    .io_in_kv(local_pes_11_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_12_io_in_inv_sum),
    .io_in_stage(local_pes_11_12_io_in_stage),
    .io_out_q(local_pes_11_12_io_out_q),
    .io_out_sum(local_pes_11_12_io_out_sum),
    .io_out_sum_exp(local_pes_11_12_io_out_sum_exp),
    .io_out_kv(local_pes_11_12_io_out_kv),
    .io_out_stage(local_pes_11_12_io_out_stage)
  );
  PE_1 local_pes_11_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_13_clock),
    .reset(local_pes_11_13_reset),
    .io_in_q(local_pes_11_13_io_in_q),
    .io_in_sum(local_pes_11_13_io_in_sum),
    .io_in_sum_exp(local_pes_11_13_io_in_sum_exp),
    .io_in_kv(local_pes_11_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_13_io_in_inv_sum),
    .io_in_stage(local_pes_11_13_io_in_stage),
    .io_out_q(local_pes_11_13_io_out_q),
    .io_out_sum(local_pes_11_13_io_out_sum),
    .io_out_sum_exp(local_pes_11_13_io_out_sum_exp),
    .io_out_kv(local_pes_11_13_io_out_kv),
    .io_out_stage(local_pes_11_13_io_out_stage)
  );
  PE_1 local_pes_11_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_14_clock),
    .reset(local_pes_11_14_reset),
    .io_in_q(local_pes_11_14_io_in_q),
    .io_in_sum(local_pes_11_14_io_in_sum),
    .io_in_sum_exp(local_pes_11_14_io_in_sum_exp),
    .io_in_kv(local_pes_11_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_14_io_in_inv_sum),
    .io_in_stage(local_pes_11_14_io_in_stage),
    .io_out_q(local_pes_11_14_io_out_q),
    .io_out_sum(local_pes_11_14_io_out_sum),
    .io_out_sum_exp(local_pes_11_14_io_out_sum_exp),
    .io_out_kv(local_pes_11_14_io_out_kv),
    .io_out_stage(local_pes_11_14_io_out_stage)
  );
  PE_1 local_pes_11_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_15_clock),
    .reset(local_pes_11_15_reset),
    .io_in_q(local_pes_11_15_io_in_q),
    .io_in_sum(local_pes_11_15_io_in_sum),
    .io_in_sum_exp(local_pes_11_15_io_in_sum_exp),
    .io_in_kv(local_pes_11_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_15_io_in_inv_sum),
    .io_in_stage(local_pes_11_15_io_in_stage),
    .io_out_q(local_pes_11_15_io_out_q),
    .io_out_sum(local_pes_11_15_io_out_sum),
    .io_out_sum_exp(local_pes_11_15_io_out_sum_exp),
    .io_out_kv(local_pes_11_15_io_out_kv),
    .io_out_stage(local_pes_11_15_io_out_stage)
  );
  PE_1 local_pes_11_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_16_clock),
    .reset(local_pes_11_16_reset),
    .io_in_q(local_pes_11_16_io_in_q),
    .io_in_sum(local_pes_11_16_io_in_sum),
    .io_in_sum_exp(local_pes_11_16_io_in_sum_exp),
    .io_in_kv(local_pes_11_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_16_io_in_inv_sum),
    .io_in_stage(local_pes_11_16_io_in_stage),
    .io_out_q(local_pes_11_16_io_out_q),
    .io_out_sum(local_pes_11_16_io_out_sum),
    .io_out_sum_exp(local_pes_11_16_io_out_sum_exp),
    .io_out_kv(local_pes_11_16_io_out_kv),
    .io_out_stage(local_pes_11_16_io_out_stage)
  );
  PE_1 local_pes_11_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_17_clock),
    .reset(local_pes_11_17_reset),
    .io_in_q(local_pes_11_17_io_in_q),
    .io_in_sum(local_pes_11_17_io_in_sum),
    .io_in_sum_exp(local_pes_11_17_io_in_sum_exp),
    .io_in_kv(local_pes_11_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_17_io_in_inv_sum),
    .io_in_stage(local_pes_11_17_io_in_stage),
    .io_out_q(local_pes_11_17_io_out_q),
    .io_out_sum(local_pes_11_17_io_out_sum),
    .io_out_sum_exp(local_pes_11_17_io_out_sum_exp),
    .io_out_kv(local_pes_11_17_io_out_kv),
    .io_out_stage(local_pes_11_17_io_out_stage)
  );
  PE_1 local_pes_11_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_18_clock),
    .reset(local_pes_11_18_reset),
    .io_in_q(local_pes_11_18_io_in_q),
    .io_in_sum(local_pes_11_18_io_in_sum),
    .io_in_sum_exp(local_pes_11_18_io_in_sum_exp),
    .io_in_kv(local_pes_11_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_18_io_in_inv_sum),
    .io_in_stage(local_pes_11_18_io_in_stage),
    .io_out_q(local_pes_11_18_io_out_q),
    .io_out_sum(local_pes_11_18_io_out_sum),
    .io_out_sum_exp(local_pes_11_18_io_out_sum_exp),
    .io_out_kv(local_pes_11_18_io_out_kv),
    .io_out_stage(local_pes_11_18_io_out_stage)
  );
  PE_1 local_pes_11_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_19_clock),
    .reset(local_pes_11_19_reset),
    .io_in_q(local_pes_11_19_io_in_q),
    .io_in_sum(local_pes_11_19_io_in_sum),
    .io_in_sum_exp(local_pes_11_19_io_in_sum_exp),
    .io_in_kv(local_pes_11_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_19_io_in_inv_sum),
    .io_in_stage(local_pes_11_19_io_in_stage),
    .io_out_q(local_pes_11_19_io_out_q),
    .io_out_sum(local_pes_11_19_io_out_sum),
    .io_out_sum_exp(local_pes_11_19_io_out_sum_exp),
    .io_out_kv(local_pes_11_19_io_out_kv),
    .io_out_stage(local_pes_11_19_io_out_stage)
  );
  PE_1 local_pes_11_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_20_clock),
    .reset(local_pes_11_20_reset),
    .io_in_q(local_pes_11_20_io_in_q),
    .io_in_sum(local_pes_11_20_io_in_sum),
    .io_in_sum_exp(local_pes_11_20_io_in_sum_exp),
    .io_in_kv(local_pes_11_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_20_io_in_inv_sum),
    .io_in_stage(local_pes_11_20_io_in_stage),
    .io_out_q(local_pes_11_20_io_out_q),
    .io_out_sum(local_pes_11_20_io_out_sum),
    .io_out_sum_exp(local_pes_11_20_io_out_sum_exp),
    .io_out_kv(local_pes_11_20_io_out_kv),
    .io_out_stage(local_pes_11_20_io_out_stage)
  );
  PE_1 local_pes_11_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_21_clock),
    .reset(local_pes_11_21_reset),
    .io_in_q(local_pes_11_21_io_in_q),
    .io_in_sum(local_pes_11_21_io_in_sum),
    .io_in_sum_exp(local_pes_11_21_io_in_sum_exp),
    .io_in_kv(local_pes_11_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_21_io_in_inv_sum),
    .io_in_stage(local_pes_11_21_io_in_stage),
    .io_out_q(local_pes_11_21_io_out_q),
    .io_out_sum(local_pes_11_21_io_out_sum),
    .io_out_sum_exp(local_pes_11_21_io_out_sum_exp),
    .io_out_kv(local_pes_11_21_io_out_kv),
    .io_out_stage(local_pes_11_21_io_out_stage)
  );
  PE_1 local_pes_11_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_22_clock),
    .reset(local_pes_11_22_reset),
    .io_in_q(local_pes_11_22_io_in_q),
    .io_in_sum(local_pes_11_22_io_in_sum),
    .io_in_sum_exp(local_pes_11_22_io_in_sum_exp),
    .io_in_kv(local_pes_11_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_22_io_in_inv_sum),
    .io_in_stage(local_pes_11_22_io_in_stage),
    .io_out_q(local_pes_11_22_io_out_q),
    .io_out_sum(local_pes_11_22_io_out_sum),
    .io_out_sum_exp(local_pes_11_22_io_out_sum_exp),
    .io_out_kv(local_pes_11_22_io_out_kv),
    .io_out_stage(local_pes_11_22_io_out_stage)
  );
  PE_1 local_pes_11_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_23_clock),
    .reset(local_pes_11_23_reset),
    .io_in_q(local_pes_11_23_io_in_q),
    .io_in_sum(local_pes_11_23_io_in_sum),
    .io_in_sum_exp(local_pes_11_23_io_in_sum_exp),
    .io_in_kv(local_pes_11_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_23_io_in_inv_sum),
    .io_in_stage(local_pes_11_23_io_in_stage),
    .io_out_q(local_pes_11_23_io_out_q),
    .io_out_sum(local_pes_11_23_io_out_sum),
    .io_out_sum_exp(local_pes_11_23_io_out_sum_exp),
    .io_out_kv(local_pes_11_23_io_out_kv),
    .io_out_stage(local_pes_11_23_io_out_stage)
  );
  PE_1 local_pes_11_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_24_clock),
    .reset(local_pes_11_24_reset),
    .io_in_q(local_pes_11_24_io_in_q),
    .io_in_sum(local_pes_11_24_io_in_sum),
    .io_in_sum_exp(local_pes_11_24_io_in_sum_exp),
    .io_in_kv(local_pes_11_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_24_io_in_inv_sum),
    .io_in_stage(local_pes_11_24_io_in_stage),
    .io_out_q(local_pes_11_24_io_out_q),
    .io_out_sum(local_pes_11_24_io_out_sum),
    .io_out_sum_exp(local_pes_11_24_io_out_sum_exp),
    .io_out_kv(local_pes_11_24_io_out_kv),
    .io_out_stage(local_pes_11_24_io_out_stage)
  );
  PE_1 local_pes_11_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_25_clock),
    .reset(local_pes_11_25_reset),
    .io_in_q(local_pes_11_25_io_in_q),
    .io_in_sum(local_pes_11_25_io_in_sum),
    .io_in_sum_exp(local_pes_11_25_io_in_sum_exp),
    .io_in_kv(local_pes_11_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_25_io_in_inv_sum),
    .io_in_stage(local_pes_11_25_io_in_stage),
    .io_out_q(local_pes_11_25_io_out_q),
    .io_out_sum(local_pes_11_25_io_out_sum),
    .io_out_sum_exp(local_pes_11_25_io_out_sum_exp),
    .io_out_kv(local_pes_11_25_io_out_kv),
    .io_out_stage(local_pes_11_25_io_out_stage)
  );
  PE_1 local_pes_11_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_26_clock),
    .reset(local_pes_11_26_reset),
    .io_in_q(local_pes_11_26_io_in_q),
    .io_in_sum(local_pes_11_26_io_in_sum),
    .io_in_sum_exp(local_pes_11_26_io_in_sum_exp),
    .io_in_kv(local_pes_11_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_26_io_in_inv_sum),
    .io_in_stage(local_pes_11_26_io_in_stage),
    .io_out_q(local_pes_11_26_io_out_q),
    .io_out_sum(local_pes_11_26_io_out_sum),
    .io_out_sum_exp(local_pes_11_26_io_out_sum_exp),
    .io_out_kv(local_pes_11_26_io_out_kv),
    .io_out_stage(local_pes_11_26_io_out_stage)
  );
  PE_1 local_pes_11_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_27_clock),
    .reset(local_pes_11_27_reset),
    .io_in_q(local_pes_11_27_io_in_q),
    .io_in_sum(local_pes_11_27_io_in_sum),
    .io_in_sum_exp(local_pes_11_27_io_in_sum_exp),
    .io_in_kv(local_pes_11_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_27_io_in_inv_sum),
    .io_in_stage(local_pes_11_27_io_in_stage),
    .io_out_q(local_pes_11_27_io_out_q),
    .io_out_sum(local_pes_11_27_io_out_sum),
    .io_out_sum_exp(local_pes_11_27_io_out_sum_exp),
    .io_out_kv(local_pes_11_27_io_out_kv),
    .io_out_stage(local_pes_11_27_io_out_stage)
  );
  PE_1 local_pes_11_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_28_clock),
    .reset(local_pes_11_28_reset),
    .io_in_q(local_pes_11_28_io_in_q),
    .io_in_sum(local_pes_11_28_io_in_sum),
    .io_in_sum_exp(local_pes_11_28_io_in_sum_exp),
    .io_in_kv(local_pes_11_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_28_io_in_inv_sum),
    .io_in_stage(local_pes_11_28_io_in_stage),
    .io_out_q(local_pes_11_28_io_out_q),
    .io_out_sum(local_pes_11_28_io_out_sum),
    .io_out_sum_exp(local_pes_11_28_io_out_sum_exp),
    .io_out_kv(local_pes_11_28_io_out_kv),
    .io_out_stage(local_pes_11_28_io_out_stage)
  );
  PE_1 local_pes_11_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_29_clock),
    .reset(local_pes_11_29_reset),
    .io_in_q(local_pes_11_29_io_in_q),
    .io_in_sum(local_pes_11_29_io_in_sum),
    .io_in_sum_exp(local_pes_11_29_io_in_sum_exp),
    .io_in_kv(local_pes_11_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_29_io_in_inv_sum),
    .io_in_stage(local_pes_11_29_io_in_stage),
    .io_out_q(local_pes_11_29_io_out_q),
    .io_out_sum(local_pes_11_29_io_out_sum),
    .io_out_sum_exp(local_pes_11_29_io_out_sum_exp),
    .io_out_kv(local_pes_11_29_io_out_kv),
    .io_out_stage(local_pes_11_29_io_out_stage)
  );
  PE_1 local_pes_11_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_30_clock),
    .reset(local_pes_11_30_reset),
    .io_in_q(local_pes_11_30_io_in_q),
    .io_in_sum(local_pes_11_30_io_in_sum),
    .io_in_sum_exp(local_pes_11_30_io_in_sum_exp),
    .io_in_kv(local_pes_11_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_30_io_in_inv_sum),
    .io_in_stage(local_pes_11_30_io_in_stage),
    .io_out_q(local_pes_11_30_io_out_q),
    .io_out_sum(local_pes_11_30_io_out_sum),
    .io_out_sum_exp(local_pes_11_30_io_out_sum_exp),
    .io_out_kv(local_pes_11_30_io_out_kv),
    .io_out_stage(local_pes_11_30_io_out_stage)
  );
  PE_1 local_pes_11_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_11_31_clock),
    .reset(local_pes_11_31_reset),
    .io_in_q(local_pes_11_31_io_in_q),
    .io_in_sum(local_pes_11_31_io_in_sum),
    .io_in_sum_exp(local_pes_11_31_io_in_sum_exp),
    .io_in_kv(local_pes_11_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_11_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_11_31_io_in_inv_sum),
    .io_in_stage(local_pes_11_31_io_in_stage),
    .io_out_q(local_pes_11_31_io_out_q),
    .io_out_sum(local_pes_11_31_io_out_sum),
    .io_out_sum_exp(local_pes_11_31_io_out_sum_exp),
    .io_out_kv(local_pes_11_31_io_out_kv),
    .io_out_stage(local_pes_11_31_io_out_stage)
  );
  PE local_pes_12_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_0_clock),
    .reset(local_pes_12_0_reset),
    .io_in_q(local_pes_12_0_io_in_q),
    .io_in_kv(local_pes_12_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_0_io_in_inv_sum),
    .io_in_stage(local_pes_12_0_io_in_stage),
    .io_out_q(local_pes_12_0_io_out_q),
    .io_out_sum(local_pes_12_0_io_out_sum),
    .io_out_kv(local_pes_12_0_io_out_kv),
    .io_out_stage(local_pes_12_0_io_out_stage)
  );
  PE_1 local_pes_12_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_1_clock),
    .reset(local_pes_12_1_reset),
    .io_in_q(local_pes_12_1_io_in_q),
    .io_in_sum(local_pes_12_1_io_in_sum),
    .io_in_sum_exp(local_pes_12_1_io_in_sum_exp),
    .io_in_kv(local_pes_12_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_1_io_in_inv_sum),
    .io_in_stage(local_pes_12_1_io_in_stage),
    .io_out_q(local_pes_12_1_io_out_q),
    .io_out_sum(local_pes_12_1_io_out_sum),
    .io_out_sum_exp(local_pes_12_1_io_out_sum_exp),
    .io_out_kv(local_pes_12_1_io_out_kv),
    .io_out_stage(local_pes_12_1_io_out_stage)
  );
  PE_1 local_pes_12_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_2_clock),
    .reset(local_pes_12_2_reset),
    .io_in_q(local_pes_12_2_io_in_q),
    .io_in_sum(local_pes_12_2_io_in_sum),
    .io_in_sum_exp(local_pes_12_2_io_in_sum_exp),
    .io_in_kv(local_pes_12_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_2_io_in_inv_sum),
    .io_in_stage(local_pes_12_2_io_in_stage),
    .io_out_q(local_pes_12_2_io_out_q),
    .io_out_sum(local_pes_12_2_io_out_sum),
    .io_out_sum_exp(local_pes_12_2_io_out_sum_exp),
    .io_out_kv(local_pes_12_2_io_out_kv),
    .io_out_stage(local_pes_12_2_io_out_stage)
  );
  PE_1 local_pes_12_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_3_clock),
    .reset(local_pes_12_3_reset),
    .io_in_q(local_pes_12_3_io_in_q),
    .io_in_sum(local_pes_12_3_io_in_sum),
    .io_in_sum_exp(local_pes_12_3_io_in_sum_exp),
    .io_in_kv(local_pes_12_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_3_io_in_inv_sum),
    .io_in_stage(local_pes_12_3_io_in_stage),
    .io_out_q(local_pes_12_3_io_out_q),
    .io_out_sum(local_pes_12_3_io_out_sum),
    .io_out_sum_exp(local_pes_12_3_io_out_sum_exp),
    .io_out_kv(local_pes_12_3_io_out_kv),
    .io_out_stage(local_pes_12_3_io_out_stage)
  );
  PE_1 local_pes_12_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_4_clock),
    .reset(local_pes_12_4_reset),
    .io_in_q(local_pes_12_4_io_in_q),
    .io_in_sum(local_pes_12_4_io_in_sum),
    .io_in_sum_exp(local_pes_12_4_io_in_sum_exp),
    .io_in_kv(local_pes_12_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_4_io_in_inv_sum),
    .io_in_stage(local_pes_12_4_io_in_stage),
    .io_out_q(local_pes_12_4_io_out_q),
    .io_out_sum(local_pes_12_4_io_out_sum),
    .io_out_sum_exp(local_pes_12_4_io_out_sum_exp),
    .io_out_kv(local_pes_12_4_io_out_kv),
    .io_out_stage(local_pes_12_4_io_out_stage)
  );
  PE_1 local_pes_12_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_5_clock),
    .reset(local_pes_12_5_reset),
    .io_in_q(local_pes_12_5_io_in_q),
    .io_in_sum(local_pes_12_5_io_in_sum),
    .io_in_sum_exp(local_pes_12_5_io_in_sum_exp),
    .io_in_kv(local_pes_12_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_5_io_in_inv_sum),
    .io_in_stage(local_pes_12_5_io_in_stage),
    .io_out_q(local_pes_12_5_io_out_q),
    .io_out_sum(local_pes_12_5_io_out_sum),
    .io_out_sum_exp(local_pes_12_5_io_out_sum_exp),
    .io_out_kv(local_pes_12_5_io_out_kv),
    .io_out_stage(local_pes_12_5_io_out_stage)
  );
  PE_1 local_pes_12_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_6_clock),
    .reset(local_pes_12_6_reset),
    .io_in_q(local_pes_12_6_io_in_q),
    .io_in_sum(local_pes_12_6_io_in_sum),
    .io_in_sum_exp(local_pes_12_6_io_in_sum_exp),
    .io_in_kv(local_pes_12_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_6_io_in_inv_sum),
    .io_in_stage(local_pes_12_6_io_in_stage),
    .io_out_q(local_pes_12_6_io_out_q),
    .io_out_sum(local_pes_12_6_io_out_sum),
    .io_out_sum_exp(local_pes_12_6_io_out_sum_exp),
    .io_out_kv(local_pes_12_6_io_out_kv),
    .io_out_stage(local_pes_12_6_io_out_stage)
  );
  PE_1 local_pes_12_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_7_clock),
    .reset(local_pes_12_7_reset),
    .io_in_q(local_pes_12_7_io_in_q),
    .io_in_sum(local_pes_12_7_io_in_sum),
    .io_in_sum_exp(local_pes_12_7_io_in_sum_exp),
    .io_in_kv(local_pes_12_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_7_io_in_inv_sum),
    .io_in_stage(local_pes_12_7_io_in_stage),
    .io_out_q(local_pes_12_7_io_out_q),
    .io_out_sum(local_pes_12_7_io_out_sum),
    .io_out_sum_exp(local_pes_12_7_io_out_sum_exp),
    .io_out_kv(local_pes_12_7_io_out_kv),
    .io_out_stage(local_pes_12_7_io_out_stage)
  );
  PE_1 local_pes_12_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_8_clock),
    .reset(local_pes_12_8_reset),
    .io_in_q(local_pes_12_8_io_in_q),
    .io_in_sum(local_pes_12_8_io_in_sum),
    .io_in_sum_exp(local_pes_12_8_io_in_sum_exp),
    .io_in_kv(local_pes_12_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_8_io_in_inv_sum),
    .io_in_stage(local_pes_12_8_io_in_stage),
    .io_out_q(local_pes_12_8_io_out_q),
    .io_out_sum(local_pes_12_8_io_out_sum),
    .io_out_sum_exp(local_pes_12_8_io_out_sum_exp),
    .io_out_kv(local_pes_12_8_io_out_kv),
    .io_out_stage(local_pes_12_8_io_out_stage)
  );
  PE_1 local_pes_12_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_9_clock),
    .reset(local_pes_12_9_reset),
    .io_in_q(local_pes_12_9_io_in_q),
    .io_in_sum(local_pes_12_9_io_in_sum),
    .io_in_sum_exp(local_pes_12_9_io_in_sum_exp),
    .io_in_kv(local_pes_12_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_9_io_in_inv_sum),
    .io_in_stage(local_pes_12_9_io_in_stage),
    .io_out_q(local_pes_12_9_io_out_q),
    .io_out_sum(local_pes_12_9_io_out_sum),
    .io_out_sum_exp(local_pes_12_9_io_out_sum_exp),
    .io_out_kv(local_pes_12_9_io_out_kv),
    .io_out_stage(local_pes_12_9_io_out_stage)
  );
  PE_1 local_pes_12_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_10_clock),
    .reset(local_pes_12_10_reset),
    .io_in_q(local_pes_12_10_io_in_q),
    .io_in_sum(local_pes_12_10_io_in_sum),
    .io_in_sum_exp(local_pes_12_10_io_in_sum_exp),
    .io_in_kv(local_pes_12_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_10_io_in_inv_sum),
    .io_in_stage(local_pes_12_10_io_in_stage),
    .io_out_q(local_pes_12_10_io_out_q),
    .io_out_sum(local_pes_12_10_io_out_sum),
    .io_out_sum_exp(local_pes_12_10_io_out_sum_exp),
    .io_out_kv(local_pes_12_10_io_out_kv),
    .io_out_stage(local_pes_12_10_io_out_stage)
  );
  PE_1 local_pes_12_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_11_clock),
    .reset(local_pes_12_11_reset),
    .io_in_q(local_pes_12_11_io_in_q),
    .io_in_sum(local_pes_12_11_io_in_sum),
    .io_in_sum_exp(local_pes_12_11_io_in_sum_exp),
    .io_in_kv(local_pes_12_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_11_io_in_inv_sum),
    .io_in_stage(local_pes_12_11_io_in_stage),
    .io_out_q(local_pes_12_11_io_out_q),
    .io_out_sum(local_pes_12_11_io_out_sum),
    .io_out_sum_exp(local_pes_12_11_io_out_sum_exp),
    .io_out_kv(local_pes_12_11_io_out_kv),
    .io_out_stage(local_pes_12_11_io_out_stage)
  );
  PE_1 local_pes_12_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_12_clock),
    .reset(local_pes_12_12_reset),
    .io_in_q(local_pes_12_12_io_in_q),
    .io_in_sum(local_pes_12_12_io_in_sum),
    .io_in_sum_exp(local_pes_12_12_io_in_sum_exp),
    .io_in_kv(local_pes_12_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_12_io_in_inv_sum),
    .io_in_stage(local_pes_12_12_io_in_stage),
    .io_out_q(local_pes_12_12_io_out_q),
    .io_out_sum(local_pes_12_12_io_out_sum),
    .io_out_sum_exp(local_pes_12_12_io_out_sum_exp),
    .io_out_kv(local_pes_12_12_io_out_kv),
    .io_out_stage(local_pes_12_12_io_out_stage)
  );
  PE_1 local_pes_12_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_13_clock),
    .reset(local_pes_12_13_reset),
    .io_in_q(local_pes_12_13_io_in_q),
    .io_in_sum(local_pes_12_13_io_in_sum),
    .io_in_sum_exp(local_pes_12_13_io_in_sum_exp),
    .io_in_kv(local_pes_12_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_13_io_in_inv_sum),
    .io_in_stage(local_pes_12_13_io_in_stage),
    .io_out_q(local_pes_12_13_io_out_q),
    .io_out_sum(local_pes_12_13_io_out_sum),
    .io_out_sum_exp(local_pes_12_13_io_out_sum_exp),
    .io_out_kv(local_pes_12_13_io_out_kv),
    .io_out_stage(local_pes_12_13_io_out_stage)
  );
  PE_1 local_pes_12_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_14_clock),
    .reset(local_pes_12_14_reset),
    .io_in_q(local_pes_12_14_io_in_q),
    .io_in_sum(local_pes_12_14_io_in_sum),
    .io_in_sum_exp(local_pes_12_14_io_in_sum_exp),
    .io_in_kv(local_pes_12_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_14_io_in_inv_sum),
    .io_in_stage(local_pes_12_14_io_in_stage),
    .io_out_q(local_pes_12_14_io_out_q),
    .io_out_sum(local_pes_12_14_io_out_sum),
    .io_out_sum_exp(local_pes_12_14_io_out_sum_exp),
    .io_out_kv(local_pes_12_14_io_out_kv),
    .io_out_stage(local_pes_12_14_io_out_stage)
  );
  PE_1 local_pes_12_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_15_clock),
    .reset(local_pes_12_15_reset),
    .io_in_q(local_pes_12_15_io_in_q),
    .io_in_sum(local_pes_12_15_io_in_sum),
    .io_in_sum_exp(local_pes_12_15_io_in_sum_exp),
    .io_in_kv(local_pes_12_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_15_io_in_inv_sum),
    .io_in_stage(local_pes_12_15_io_in_stage),
    .io_out_q(local_pes_12_15_io_out_q),
    .io_out_sum(local_pes_12_15_io_out_sum),
    .io_out_sum_exp(local_pes_12_15_io_out_sum_exp),
    .io_out_kv(local_pes_12_15_io_out_kv),
    .io_out_stage(local_pes_12_15_io_out_stage)
  );
  PE_1 local_pes_12_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_16_clock),
    .reset(local_pes_12_16_reset),
    .io_in_q(local_pes_12_16_io_in_q),
    .io_in_sum(local_pes_12_16_io_in_sum),
    .io_in_sum_exp(local_pes_12_16_io_in_sum_exp),
    .io_in_kv(local_pes_12_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_16_io_in_inv_sum),
    .io_in_stage(local_pes_12_16_io_in_stage),
    .io_out_q(local_pes_12_16_io_out_q),
    .io_out_sum(local_pes_12_16_io_out_sum),
    .io_out_sum_exp(local_pes_12_16_io_out_sum_exp),
    .io_out_kv(local_pes_12_16_io_out_kv),
    .io_out_stage(local_pes_12_16_io_out_stage)
  );
  PE_1 local_pes_12_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_17_clock),
    .reset(local_pes_12_17_reset),
    .io_in_q(local_pes_12_17_io_in_q),
    .io_in_sum(local_pes_12_17_io_in_sum),
    .io_in_sum_exp(local_pes_12_17_io_in_sum_exp),
    .io_in_kv(local_pes_12_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_17_io_in_inv_sum),
    .io_in_stage(local_pes_12_17_io_in_stage),
    .io_out_q(local_pes_12_17_io_out_q),
    .io_out_sum(local_pes_12_17_io_out_sum),
    .io_out_sum_exp(local_pes_12_17_io_out_sum_exp),
    .io_out_kv(local_pes_12_17_io_out_kv),
    .io_out_stage(local_pes_12_17_io_out_stage)
  );
  PE_1 local_pes_12_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_18_clock),
    .reset(local_pes_12_18_reset),
    .io_in_q(local_pes_12_18_io_in_q),
    .io_in_sum(local_pes_12_18_io_in_sum),
    .io_in_sum_exp(local_pes_12_18_io_in_sum_exp),
    .io_in_kv(local_pes_12_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_18_io_in_inv_sum),
    .io_in_stage(local_pes_12_18_io_in_stage),
    .io_out_q(local_pes_12_18_io_out_q),
    .io_out_sum(local_pes_12_18_io_out_sum),
    .io_out_sum_exp(local_pes_12_18_io_out_sum_exp),
    .io_out_kv(local_pes_12_18_io_out_kv),
    .io_out_stage(local_pes_12_18_io_out_stage)
  );
  PE_1 local_pes_12_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_19_clock),
    .reset(local_pes_12_19_reset),
    .io_in_q(local_pes_12_19_io_in_q),
    .io_in_sum(local_pes_12_19_io_in_sum),
    .io_in_sum_exp(local_pes_12_19_io_in_sum_exp),
    .io_in_kv(local_pes_12_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_19_io_in_inv_sum),
    .io_in_stage(local_pes_12_19_io_in_stage),
    .io_out_q(local_pes_12_19_io_out_q),
    .io_out_sum(local_pes_12_19_io_out_sum),
    .io_out_sum_exp(local_pes_12_19_io_out_sum_exp),
    .io_out_kv(local_pes_12_19_io_out_kv),
    .io_out_stage(local_pes_12_19_io_out_stage)
  );
  PE_1 local_pes_12_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_20_clock),
    .reset(local_pes_12_20_reset),
    .io_in_q(local_pes_12_20_io_in_q),
    .io_in_sum(local_pes_12_20_io_in_sum),
    .io_in_sum_exp(local_pes_12_20_io_in_sum_exp),
    .io_in_kv(local_pes_12_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_20_io_in_inv_sum),
    .io_in_stage(local_pes_12_20_io_in_stage),
    .io_out_q(local_pes_12_20_io_out_q),
    .io_out_sum(local_pes_12_20_io_out_sum),
    .io_out_sum_exp(local_pes_12_20_io_out_sum_exp),
    .io_out_kv(local_pes_12_20_io_out_kv),
    .io_out_stage(local_pes_12_20_io_out_stage)
  );
  PE_1 local_pes_12_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_21_clock),
    .reset(local_pes_12_21_reset),
    .io_in_q(local_pes_12_21_io_in_q),
    .io_in_sum(local_pes_12_21_io_in_sum),
    .io_in_sum_exp(local_pes_12_21_io_in_sum_exp),
    .io_in_kv(local_pes_12_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_21_io_in_inv_sum),
    .io_in_stage(local_pes_12_21_io_in_stage),
    .io_out_q(local_pes_12_21_io_out_q),
    .io_out_sum(local_pes_12_21_io_out_sum),
    .io_out_sum_exp(local_pes_12_21_io_out_sum_exp),
    .io_out_kv(local_pes_12_21_io_out_kv),
    .io_out_stage(local_pes_12_21_io_out_stage)
  );
  PE_1 local_pes_12_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_22_clock),
    .reset(local_pes_12_22_reset),
    .io_in_q(local_pes_12_22_io_in_q),
    .io_in_sum(local_pes_12_22_io_in_sum),
    .io_in_sum_exp(local_pes_12_22_io_in_sum_exp),
    .io_in_kv(local_pes_12_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_22_io_in_inv_sum),
    .io_in_stage(local_pes_12_22_io_in_stage),
    .io_out_q(local_pes_12_22_io_out_q),
    .io_out_sum(local_pes_12_22_io_out_sum),
    .io_out_sum_exp(local_pes_12_22_io_out_sum_exp),
    .io_out_kv(local_pes_12_22_io_out_kv),
    .io_out_stage(local_pes_12_22_io_out_stage)
  );
  PE_1 local_pes_12_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_23_clock),
    .reset(local_pes_12_23_reset),
    .io_in_q(local_pes_12_23_io_in_q),
    .io_in_sum(local_pes_12_23_io_in_sum),
    .io_in_sum_exp(local_pes_12_23_io_in_sum_exp),
    .io_in_kv(local_pes_12_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_23_io_in_inv_sum),
    .io_in_stage(local_pes_12_23_io_in_stage),
    .io_out_q(local_pes_12_23_io_out_q),
    .io_out_sum(local_pes_12_23_io_out_sum),
    .io_out_sum_exp(local_pes_12_23_io_out_sum_exp),
    .io_out_kv(local_pes_12_23_io_out_kv),
    .io_out_stage(local_pes_12_23_io_out_stage)
  );
  PE_1 local_pes_12_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_24_clock),
    .reset(local_pes_12_24_reset),
    .io_in_q(local_pes_12_24_io_in_q),
    .io_in_sum(local_pes_12_24_io_in_sum),
    .io_in_sum_exp(local_pes_12_24_io_in_sum_exp),
    .io_in_kv(local_pes_12_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_24_io_in_inv_sum),
    .io_in_stage(local_pes_12_24_io_in_stage),
    .io_out_q(local_pes_12_24_io_out_q),
    .io_out_sum(local_pes_12_24_io_out_sum),
    .io_out_sum_exp(local_pes_12_24_io_out_sum_exp),
    .io_out_kv(local_pes_12_24_io_out_kv),
    .io_out_stage(local_pes_12_24_io_out_stage)
  );
  PE_1 local_pes_12_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_25_clock),
    .reset(local_pes_12_25_reset),
    .io_in_q(local_pes_12_25_io_in_q),
    .io_in_sum(local_pes_12_25_io_in_sum),
    .io_in_sum_exp(local_pes_12_25_io_in_sum_exp),
    .io_in_kv(local_pes_12_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_25_io_in_inv_sum),
    .io_in_stage(local_pes_12_25_io_in_stage),
    .io_out_q(local_pes_12_25_io_out_q),
    .io_out_sum(local_pes_12_25_io_out_sum),
    .io_out_sum_exp(local_pes_12_25_io_out_sum_exp),
    .io_out_kv(local_pes_12_25_io_out_kv),
    .io_out_stage(local_pes_12_25_io_out_stage)
  );
  PE_1 local_pes_12_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_26_clock),
    .reset(local_pes_12_26_reset),
    .io_in_q(local_pes_12_26_io_in_q),
    .io_in_sum(local_pes_12_26_io_in_sum),
    .io_in_sum_exp(local_pes_12_26_io_in_sum_exp),
    .io_in_kv(local_pes_12_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_26_io_in_inv_sum),
    .io_in_stage(local_pes_12_26_io_in_stage),
    .io_out_q(local_pes_12_26_io_out_q),
    .io_out_sum(local_pes_12_26_io_out_sum),
    .io_out_sum_exp(local_pes_12_26_io_out_sum_exp),
    .io_out_kv(local_pes_12_26_io_out_kv),
    .io_out_stage(local_pes_12_26_io_out_stage)
  );
  PE_1 local_pes_12_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_27_clock),
    .reset(local_pes_12_27_reset),
    .io_in_q(local_pes_12_27_io_in_q),
    .io_in_sum(local_pes_12_27_io_in_sum),
    .io_in_sum_exp(local_pes_12_27_io_in_sum_exp),
    .io_in_kv(local_pes_12_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_27_io_in_inv_sum),
    .io_in_stage(local_pes_12_27_io_in_stage),
    .io_out_q(local_pes_12_27_io_out_q),
    .io_out_sum(local_pes_12_27_io_out_sum),
    .io_out_sum_exp(local_pes_12_27_io_out_sum_exp),
    .io_out_kv(local_pes_12_27_io_out_kv),
    .io_out_stage(local_pes_12_27_io_out_stage)
  );
  PE_1 local_pes_12_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_28_clock),
    .reset(local_pes_12_28_reset),
    .io_in_q(local_pes_12_28_io_in_q),
    .io_in_sum(local_pes_12_28_io_in_sum),
    .io_in_sum_exp(local_pes_12_28_io_in_sum_exp),
    .io_in_kv(local_pes_12_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_28_io_in_inv_sum),
    .io_in_stage(local_pes_12_28_io_in_stage),
    .io_out_q(local_pes_12_28_io_out_q),
    .io_out_sum(local_pes_12_28_io_out_sum),
    .io_out_sum_exp(local_pes_12_28_io_out_sum_exp),
    .io_out_kv(local_pes_12_28_io_out_kv),
    .io_out_stage(local_pes_12_28_io_out_stage)
  );
  PE_1 local_pes_12_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_29_clock),
    .reset(local_pes_12_29_reset),
    .io_in_q(local_pes_12_29_io_in_q),
    .io_in_sum(local_pes_12_29_io_in_sum),
    .io_in_sum_exp(local_pes_12_29_io_in_sum_exp),
    .io_in_kv(local_pes_12_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_29_io_in_inv_sum),
    .io_in_stage(local_pes_12_29_io_in_stage),
    .io_out_q(local_pes_12_29_io_out_q),
    .io_out_sum(local_pes_12_29_io_out_sum),
    .io_out_sum_exp(local_pes_12_29_io_out_sum_exp),
    .io_out_kv(local_pes_12_29_io_out_kv),
    .io_out_stage(local_pes_12_29_io_out_stage)
  );
  PE_1 local_pes_12_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_30_clock),
    .reset(local_pes_12_30_reset),
    .io_in_q(local_pes_12_30_io_in_q),
    .io_in_sum(local_pes_12_30_io_in_sum),
    .io_in_sum_exp(local_pes_12_30_io_in_sum_exp),
    .io_in_kv(local_pes_12_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_30_io_in_inv_sum),
    .io_in_stage(local_pes_12_30_io_in_stage),
    .io_out_q(local_pes_12_30_io_out_q),
    .io_out_sum(local_pes_12_30_io_out_sum),
    .io_out_sum_exp(local_pes_12_30_io_out_sum_exp),
    .io_out_kv(local_pes_12_30_io_out_kv),
    .io_out_stage(local_pes_12_30_io_out_stage)
  );
  PE_1 local_pes_12_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_12_31_clock),
    .reset(local_pes_12_31_reset),
    .io_in_q(local_pes_12_31_io_in_q),
    .io_in_sum(local_pes_12_31_io_in_sum),
    .io_in_sum_exp(local_pes_12_31_io_in_sum_exp),
    .io_in_kv(local_pes_12_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_12_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_12_31_io_in_inv_sum),
    .io_in_stage(local_pes_12_31_io_in_stage),
    .io_out_q(local_pes_12_31_io_out_q),
    .io_out_sum(local_pes_12_31_io_out_sum),
    .io_out_sum_exp(local_pes_12_31_io_out_sum_exp),
    .io_out_kv(local_pes_12_31_io_out_kv),
    .io_out_stage(local_pes_12_31_io_out_stage)
  );
  PE local_pes_13_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_0_clock),
    .reset(local_pes_13_0_reset),
    .io_in_q(local_pes_13_0_io_in_q),
    .io_in_kv(local_pes_13_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_0_io_in_inv_sum),
    .io_in_stage(local_pes_13_0_io_in_stage),
    .io_out_q(local_pes_13_0_io_out_q),
    .io_out_sum(local_pes_13_0_io_out_sum),
    .io_out_kv(local_pes_13_0_io_out_kv),
    .io_out_stage(local_pes_13_0_io_out_stage)
  );
  PE_1 local_pes_13_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_1_clock),
    .reset(local_pes_13_1_reset),
    .io_in_q(local_pes_13_1_io_in_q),
    .io_in_sum(local_pes_13_1_io_in_sum),
    .io_in_sum_exp(local_pes_13_1_io_in_sum_exp),
    .io_in_kv(local_pes_13_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_1_io_in_inv_sum),
    .io_in_stage(local_pes_13_1_io_in_stage),
    .io_out_q(local_pes_13_1_io_out_q),
    .io_out_sum(local_pes_13_1_io_out_sum),
    .io_out_sum_exp(local_pes_13_1_io_out_sum_exp),
    .io_out_kv(local_pes_13_1_io_out_kv),
    .io_out_stage(local_pes_13_1_io_out_stage)
  );
  PE_1 local_pes_13_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_2_clock),
    .reset(local_pes_13_2_reset),
    .io_in_q(local_pes_13_2_io_in_q),
    .io_in_sum(local_pes_13_2_io_in_sum),
    .io_in_sum_exp(local_pes_13_2_io_in_sum_exp),
    .io_in_kv(local_pes_13_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_2_io_in_inv_sum),
    .io_in_stage(local_pes_13_2_io_in_stage),
    .io_out_q(local_pes_13_2_io_out_q),
    .io_out_sum(local_pes_13_2_io_out_sum),
    .io_out_sum_exp(local_pes_13_2_io_out_sum_exp),
    .io_out_kv(local_pes_13_2_io_out_kv),
    .io_out_stage(local_pes_13_2_io_out_stage)
  );
  PE_1 local_pes_13_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_3_clock),
    .reset(local_pes_13_3_reset),
    .io_in_q(local_pes_13_3_io_in_q),
    .io_in_sum(local_pes_13_3_io_in_sum),
    .io_in_sum_exp(local_pes_13_3_io_in_sum_exp),
    .io_in_kv(local_pes_13_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_3_io_in_inv_sum),
    .io_in_stage(local_pes_13_3_io_in_stage),
    .io_out_q(local_pes_13_3_io_out_q),
    .io_out_sum(local_pes_13_3_io_out_sum),
    .io_out_sum_exp(local_pes_13_3_io_out_sum_exp),
    .io_out_kv(local_pes_13_3_io_out_kv),
    .io_out_stage(local_pes_13_3_io_out_stage)
  );
  PE_1 local_pes_13_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_4_clock),
    .reset(local_pes_13_4_reset),
    .io_in_q(local_pes_13_4_io_in_q),
    .io_in_sum(local_pes_13_4_io_in_sum),
    .io_in_sum_exp(local_pes_13_4_io_in_sum_exp),
    .io_in_kv(local_pes_13_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_4_io_in_inv_sum),
    .io_in_stage(local_pes_13_4_io_in_stage),
    .io_out_q(local_pes_13_4_io_out_q),
    .io_out_sum(local_pes_13_4_io_out_sum),
    .io_out_sum_exp(local_pes_13_4_io_out_sum_exp),
    .io_out_kv(local_pes_13_4_io_out_kv),
    .io_out_stage(local_pes_13_4_io_out_stage)
  );
  PE_1 local_pes_13_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_5_clock),
    .reset(local_pes_13_5_reset),
    .io_in_q(local_pes_13_5_io_in_q),
    .io_in_sum(local_pes_13_5_io_in_sum),
    .io_in_sum_exp(local_pes_13_5_io_in_sum_exp),
    .io_in_kv(local_pes_13_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_5_io_in_inv_sum),
    .io_in_stage(local_pes_13_5_io_in_stage),
    .io_out_q(local_pes_13_5_io_out_q),
    .io_out_sum(local_pes_13_5_io_out_sum),
    .io_out_sum_exp(local_pes_13_5_io_out_sum_exp),
    .io_out_kv(local_pes_13_5_io_out_kv),
    .io_out_stage(local_pes_13_5_io_out_stage)
  );
  PE_1 local_pes_13_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_6_clock),
    .reset(local_pes_13_6_reset),
    .io_in_q(local_pes_13_6_io_in_q),
    .io_in_sum(local_pes_13_6_io_in_sum),
    .io_in_sum_exp(local_pes_13_6_io_in_sum_exp),
    .io_in_kv(local_pes_13_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_6_io_in_inv_sum),
    .io_in_stage(local_pes_13_6_io_in_stage),
    .io_out_q(local_pes_13_6_io_out_q),
    .io_out_sum(local_pes_13_6_io_out_sum),
    .io_out_sum_exp(local_pes_13_6_io_out_sum_exp),
    .io_out_kv(local_pes_13_6_io_out_kv),
    .io_out_stage(local_pes_13_6_io_out_stage)
  );
  PE_1 local_pes_13_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_7_clock),
    .reset(local_pes_13_7_reset),
    .io_in_q(local_pes_13_7_io_in_q),
    .io_in_sum(local_pes_13_7_io_in_sum),
    .io_in_sum_exp(local_pes_13_7_io_in_sum_exp),
    .io_in_kv(local_pes_13_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_7_io_in_inv_sum),
    .io_in_stage(local_pes_13_7_io_in_stage),
    .io_out_q(local_pes_13_7_io_out_q),
    .io_out_sum(local_pes_13_7_io_out_sum),
    .io_out_sum_exp(local_pes_13_7_io_out_sum_exp),
    .io_out_kv(local_pes_13_7_io_out_kv),
    .io_out_stage(local_pes_13_7_io_out_stage)
  );
  PE_1 local_pes_13_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_8_clock),
    .reset(local_pes_13_8_reset),
    .io_in_q(local_pes_13_8_io_in_q),
    .io_in_sum(local_pes_13_8_io_in_sum),
    .io_in_sum_exp(local_pes_13_8_io_in_sum_exp),
    .io_in_kv(local_pes_13_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_8_io_in_inv_sum),
    .io_in_stage(local_pes_13_8_io_in_stage),
    .io_out_q(local_pes_13_8_io_out_q),
    .io_out_sum(local_pes_13_8_io_out_sum),
    .io_out_sum_exp(local_pes_13_8_io_out_sum_exp),
    .io_out_kv(local_pes_13_8_io_out_kv),
    .io_out_stage(local_pes_13_8_io_out_stage)
  );
  PE_1 local_pes_13_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_9_clock),
    .reset(local_pes_13_9_reset),
    .io_in_q(local_pes_13_9_io_in_q),
    .io_in_sum(local_pes_13_9_io_in_sum),
    .io_in_sum_exp(local_pes_13_9_io_in_sum_exp),
    .io_in_kv(local_pes_13_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_9_io_in_inv_sum),
    .io_in_stage(local_pes_13_9_io_in_stage),
    .io_out_q(local_pes_13_9_io_out_q),
    .io_out_sum(local_pes_13_9_io_out_sum),
    .io_out_sum_exp(local_pes_13_9_io_out_sum_exp),
    .io_out_kv(local_pes_13_9_io_out_kv),
    .io_out_stage(local_pes_13_9_io_out_stage)
  );
  PE_1 local_pes_13_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_10_clock),
    .reset(local_pes_13_10_reset),
    .io_in_q(local_pes_13_10_io_in_q),
    .io_in_sum(local_pes_13_10_io_in_sum),
    .io_in_sum_exp(local_pes_13_10_io_in_sum_exp),
    .io_in_kv(local_pes_13_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_10_io_in_inv_sum),
    .io_in_stage(local_pes_13_10_io_in_stage),
    .io_out_q(local_pes_13_10_io_out_q),
    .io_out_sum(local_pes_13_10_io_out_sum),
    .io_out_sum_exp(local_pes_13_10_io_out_sum_exp),
    .io_out_kv(local_pes_13_10_io_out_kv),
    .io_out_stage(local_pes_13_10_io_out_stage)
  );
  PE_1 local_pes_13_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_11_clock),
    .reset(local_pes_13_11_reset),
    .io_in_q(local_pes_13_11_io_in_q),
    .io_in_sum(local_pes_13_11_io_in_sum),
    .io_in_sum_exp(local_pes_13_11_io_in_sum_exp),
    .io_in_kv(local_pes_13_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_11_io_in_inv_sum),
    .io_in_stage(local_pes_13_11_io_in_stage),
    .io_out_q(local_pes_13_11_io_out_q),
    .io_out_sum(local_pes_13_11_io_out_sum),
    .io_out_sum_exp(local_pes_13_11_io_out_sum_exp),
    .io_out_kv(local_pes_13_11_io_out_kv),
    .io_out_stage(local_pes_13_11_io_out_stage)
  );
  PE_1 local_pes_13_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_12_clock),
    .reset(local_pes_13_12_reset),
    .io_in_q(local_pes_13_12_io_in_q),
    .io_in_sum(local_pes_13_12_io_in_sum),
    .io_in_sum_exp(local_pes_13_12_io_in_sum_exp),
    .io_in_kv(local_pes_13_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_12_io_in_inv_sum),
    .io_in_stage(local_pes_13_12_io_in_stage),
    .io_out_q(local_pes_13_12_io_out_q),
    .io_out_sum(local_pes_13_12_io_out_sum),
    .io_out_sum_exp(local_pes_13_12_io_out_sum_exp),
    .io_out_kv(local_pes_13_12_io_out_kv),
    .io_out_stage(local_pes_13_12_io_out_stage)
  );
  PE_1 local_pes_13_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_13_clock),
    .reset(local_pes_13_13_reset),
    .io_in_q(local_pes_13_13_io_in_q),
    .io_in_sum(local_pes_13_13_io_in_sum),
    .io_in_sum_exp(local_pes_13_13_io_in_sum_exp),
    .io_in_kv(local_pes_13_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_13_io_in_inv_sum),
    .io_in_stage(local_pes_13_13_io_in_stage),
    .io_out_q(local_pes_13_13_io_out_q),
    .io_out_sum(local_pes_13_13_io_out_sum),
    .io_out_sum_exp(local_pes_13_13_io_out_sum_exp),
    .io_out_kv(local_pes_13_13_io_out_kv),
    .io_out_stage(local_pes_13_13_io_out_stage)
  );
  PE_1 local_pes_13_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_14_clock),
    .reset(local_pes_13_14_reset),
    .io_in_q(local_pes_13_14_io_in_q),
    .io_in_sum(local_pes_13_14_io_in_sum),
    .io_in_sum_exp(local_pes_13_14_io_in_sum_exp),
    .io_in_kv(local_pes_13_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_14_io_in_inv_sum),
    .io_in_stage(local_pes_13_14_io_in_stage),
    .io_out_q(local_pes_13_14_io_out_q),
    .io_out_sum(local_pes_13_14_io_out_sum),
    .io_out_sum_exp(local_pes_13_14_io_out_sum_exp),
    .io_out_kv(local_pes_13_14_io_out_kv),
    .io_out_stage(local_pes_13_14_io_out_stage)
  );
  PE_1 local_pes_13_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_15_clock),
    .reset(local_pes_13_15_reset),
    .io_in_q(local_pes_13_15_io_in_q),
    .io_in_sum(local_pes_13_15_io_in_sum),
    .io_in_sum_exp(local_pes_13_15_io_in_sum_exp),
    .io_in_kv(local_pes_13_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_15_io_in_inv_sum),
    .io_in_stage(local_pes_13_15_io_in_stage),
    .io_out_q(local_pes_13_15_io_out_q),
    .io_out_sum(local_pes_13_15_io_out_sum),
    .io_out_sum_exp(local_pes_13_15_io_out_sum_exp),
    .io_out_kv(local_pes_13_15_io_out_kv),
    .io_out_stage(local_pes_13_15_io_out_stage)
  );
  PE_1 local_pes_13_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_16_clock),
    .reset(local_pes_13_16_reset),
    .io_in_q(local_pes_13_16_io_in_q),
    .io_in_sum(local_pes_13_16_io_in_sum),
    .io_in_sum_exp(local_pes_13_16_io_in_sum_exp),
    .io_in_kv(local_pes_13_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_16_io_in_inv_sum),
    .io_in_stage(local_pes_13_16_io_in_stage),
    .io_out_q(local_pes_13_16_io_out_q),
    .io_out_sum(local_pes_13_16_io_out_sum),
    .io_out_sum_exp(local_pes_13_16_io_out_sum_exp),
    .io_out_kv(local_pes_13_16_io_out_kv),
    .io_out_stage(local_pes_13_16_io_out_stage)
  );
  PE_1 local_pes_13_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_17_clock),
    .reset(local_pes_13_17_reset),
    .io_in_q(local_pes_13_17_io_in_q),
    .io_in_sum(local_pes_13_17_io_in_sum),
    .io_in_sum_exp(local_pes_13_17_io_in_sum_exp),
    .io_in_kv(local_pes_13_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_17_io_in_inv_sum),
    .io_in_stage(local_pes_13_17_io_in_stage),
    .io_out_q(local_pes_13_17_io_out_q),
    .io_out_sum(local_pes_13_17_io_out_sum),
    .io_out_sum_exp(local_pes_13_17_io_out_sum_exp),
    .io_out_kv(local_pes_13_17_io_out_kv),
    .io_out_stage(local_pes_13_17_io_out_stage)
  );
  PE_1 local_pes_13_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_18_clock),
    .reset(local_pes_13_18_reset),
    .io_in_q(local_pes_13_18_io_in_q),
    .io_in_sum(local_pes_13_18_io_in_sum),
    .io_in_sum_exp(local_pes_13_18_io_in_sum_exp),
    .io_in_kv(local_pes_13_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_18_io_in_inv_sum),
    .io_in_stage(local_pes_13_18_io_in_stage),
    .io_out_q(local_pes_13_18_io_out_q),
    .io_out_sum(local_pes_13_18_io_out_sum),
    .io_out_sum_exp(local_pes_13_18_io_out_sum_exp),
    .io_out_kv(local_pes_13_18_io_out_kv),
    .io_out_stage(local_pes_13_18_io_out_stage)
  );
  PE_1 local_pes_13_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_19_clock),
    .reset(local_pes_13_19_reset),
    .io_in_q(local_pes_13_19_io_in_q),
    .io_in_sum(local_pes_13_19_io_in_sum),
    .io_in_sum_exp(local_pes_13_19_io_in_sum_exp),
    .io_in_kv(local_pes_13_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_19_io_in_inv_sum),
    .io_in_stage(local_pes_13_19_io_in_stage),
    .io_out_q(local_pes_13_19_io_out_q),
    .io_out_sum(local_pes_13_19_io_out_sum),
    .io_out_sum_exp(local_pes_13_19_io_out_sum_exp),
    .io_out_kv(local_pes_13_19_io_out_kv),
    .io_out_stage(local_pes_13_19_io_out_stage)
  );
  PE_1 local_pes_13_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_20_clock),
    .reset(local_pes_13_20_reset),
    .io_in_q(local_pes_13_20_io_in_q),
    .io_in_sum(local_pes_13_20_io_in_sum),
    .io_in_sum_exp(local_pes_13_20_io_in_sum_exp),
    .io_in_kv(local_pes_13_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_20_io_in_inv_sum),
    .io_in_stage(local_pes_13_20_io_in_stage),
    .io_out_q(local_pes_13_20_io_out_q),
    .io_out_sum(local_pes_13_20_io_out_sum),
    .io_out_sum_exp(local_pes_13_20_io_out_sum_exp),
    .io_out_kv(local_pes_13_20_io_out_kv),
    .io_out_stage(local_pes_13_20_io_out_stage)
  );
  PE_1 local_pes_13_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_21_clock),
    .reset(local_pes_13_21_reset),
    .io_in_q(local_pes_13_21_io_in_q),
    .io_in_sum(local_pes_13_21_io_in_sum),
    .io_in_sum_exp(local_pes_13_21_io_in_sum_exp),
    .io_in_kv(local_pes_13_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_21_io_in_inv_sum),
    .io_in_stage(local_pes_13_21_io_in_stage),
    .io_out_q(local_pes_13_21_io_out_q),
    .io_out_sum(local_pes_13_21_io_out_sum),
    .io_out_sum_exp(local_pes_13_21_io_out_sum_exp),
    .io_out_kv(local_pes_13_21_io_out_kv),
    .io_out_stage(local_pes_13_21_io_out_stage)
  );
  PE_1 local_pes_13_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_22_clock),
    .reset(local_pes_13_22_reset),
    .io_in_q(local_pes_13_22_io_in_q),
    .io_in_sum(local_pes_13_22_io_in_sum),
    .io_in_sum_exp(local_pes_13_22_io_in_sum_exp),
    .io_in_kv(local_pes_13_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_22_io_in_inv_sum),
    .io_in_stage(local_pes_13_22_io_in_stage),
    .io_out_q(local_pes_13_22_io_out_q),
    .io_out_sum(local_pes_13_22_io_out_sum),
    .io_out_sum_exp(local_pes_13_22_io_out_sum_exp),
    .io_out_kv(local_pes_13_22_io_out_kv),
    .io_out_stage(local_pes_13_22_io_out_stage)
  );
  PE_1 local_pes_13_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_23_clock),
    .reset(local_pes_13_23_reset),
    .io_in_q(local_pes_13_23_io_in_q),
    .io_in_sum(local_pes_13_23_io_in_sum),
    .io_in_sum_exp(local_pes_13_23_io_in_sum_exp),
    .io_in_kv(local_pes_13_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_23_io_in_inv_sum),
    .io_in_stage(local_pes_13_23_io_in_stage),
    .io_out_q(local_pes_13_23_io_out_q),
    .io_out_sum(local_pes_13_23_io_out_sum),
    .io_out_sum_exp(local_pes_13_23_io_out_sum_exp),
    .io_out_kv(local_pes_13_23_io_out_kv),
    .io_out_stage(local_pes_13_23_io_out_stage)
  );
  PE_1 local_pes_13_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_24_clock),
    .reset(local_pes_13_24_reset),
    .io_in_q(local_pes_13_24_io_in_q),
    .io_in_sum(local_pes_13_24_io_in_sum),
    .io_in_sum_exp(local_pes_13_24_io_in_sum_exp),
    .io_in_kv(local_pes_13_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_24_io_in_inv_sum),
    .io_in_stage(local_pes_13_24_io_in_stage),
    .io_out_q(local_pes_13_24_io_out_q),
    .io_out_sum(local_pes_13_24_io_out_sum),
    .io_out_sum_exp(local_pes_13_24_io_out_sum_exp),
    .io_out_kv(local_pes_13_24_io_out_kv),
    .io_out_stage(local_pes_13_24_io_out_stage)
  );
  PE_1 local_pes_13_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_25_clock),
    .reset(local_pes_13_25_reset),
    .io_in_q(local_pes_13_25_io_in_q),
    .io_in_sum(local_pes_13_25_io_in_sum),
    .io_in_sum_exp(local_pes_13_25_io_in_sum_exp),
    .io_in_kv(local_pes_13_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_25_io_in_inv_sum),
    .io_in_stage(local_pes_13_25_io_in_stage),
    .io_out_q(local_pes_13_25_io_out_q),
    .io_out_sum(local_pes_13_25_io_out_sum),
    .io_out_sum_exp(local_pes_13_25_io_out_sum_exp),
    .io_out_kv(local_pes_13_25_io_out_kv),
    .io_out_stage(local_pes_13_25_io_out_stage)
  );
  PE_1 local_pes_13_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_26_clock),
    .reset(local_pes_13_26_reset),
    .io_in_q(local_pes_13_26_io_in_q),
    .io_in_sum(local_pes_13_26_io_in_sum),
    .io_in_sum_exp(local_pes_13_26_io_in_sum_exp),
    .io_in_kv(local_pes_13_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_26_io_in_inv_sum),
    .io_in_stage(local_pes_13_26_io_in_stage),
    .io_out_q(local_pes_13_26_io_out_q),
    .io_out_sum(local_pes_13_26_io_out_sum),
    .io_out_sum_exp(local_pes_13_26_io_out_sum_exp),
    .io_out_kv(local_pes_13_26_io_out_kv),
    .io_out_stage(local_pes_13_26_io_out_stage)
  );
  PE_1 local_pes_13_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_27_clock),
    .reset(local_pes_13_27_reset),
    .io_in_q(local_pes_13_27_io_in_q),
    .io_in_sum(local_pes_13_27_io_in_sum),
    .io_in_sum_exp(local_pes_13_27_io_in_sum_exp),
    .io_in_kv(local_pes_13_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_27_io_in_inv_sum),
    .io_in_stage(local_pes_13_27_io_in_stage),
    .io_out_q(local_pes_13_27_io_out_q),
    .io_out_sum(local_pes_13_27_io_out_sum),
    .io_out_sum_exp(local_pes_13_27_io_out_sum_exp),
    .io_out_kv(local_pes_13_27_io_out_kv),
    .io_out_stage(local_pes_13_27_io_out_stage)
  );
  PE_1 local_pes_13_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_28_clock),
    .reset(local_pes_13_28_reset),
    .io_in_q(local_pes_13_28_io_in_q),
    .io_in_sum(local_pes_13_28_io_in_sum),
    .io_in_sum_exp(local_pes_13_28_io_in_sum_exp),
    .io_in_kv(local_pes_13_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_28_io_in_inv_sum),
    .io_in_stage(local_pes_13_28_io_in_stage),
    .io_out_q(local_pes_13_28_io_out_q),
    .io_out_sum(local_pes_13_28_io_out_sum),
    .io_out_sum_exp(local_pes_13_28_io_out_sum_exp),
    .io_out_kv(local_pes_13_28_io_out_kv),
    .io_out_stage(local_pes_13_28_io_out_stage)
  );
  PE_1 local_pes_13_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_29_clock),
    .reset(local_pes_13_29_reset),
    .io_in_q(local_pes_13_29_io_in_q),
    .io_in_sum(local_pes_13_29_io_in_sum),
    .io_in_sum_exp(local_pes_13_29_io_in_sum_exp),
    .io_in_kv(local_pes_13_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_29_io_in_inv_sum),
    .io_in_stage(local_pes_13_29_io_in_stage),
    .io_out_q(local_pes_13_29_io_out_q),
    .io_out_sum(local_pes_13_29_io_out_sum),
    .io_out_sum_exp(local_pes_13_29_io_out_sum_exp),
    .io_out_kv(local_pes_13_29_io_out_kv),
    .io_out_stage(local_pes_13_29_io_out_stage)
  );
  PE_1 local_pes_13_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_30_clock),
    .reset(local_pes_13_30_reset),
    .io_in_q(local_pes_13_30_io_in_q),
    .io_in_sum(local_pes_13_30_io_in_sum),
    .io_in_sum_exp(local_pes_13_30_io_in_sum_exp),
    .io_in_kv(local_pes_13_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_30_io_in_inv_sum),
    .io_in_stage(local_pes_13_30_io_in_stage),
    .io_out_q(local_pes_13_30_io_out_q),
    .io_out_sum(local_pes_13_30_io_out_sum),
    .io_out_sum_exp(local_pes_13_30_io_out_sum_exp),
    .io_out_kv(local_pes_13_30_io_out_kv),
    .io_out_stage(local_pes_13_30_io_out_stage)
  );
  PE_1 local_pes_13_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_13_31_clock),
    .reset(local_pes_13_31_reset),
    .io_in_q(local_pes_13_31_io_in_q),
    .io_in_sum(local_pes_13_31_io_in_sum),
    .io_in_sum_exp(local_pes_13_31_io_in_sum_exp),
    .io_in_kv(local_pes_13_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_13_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_13_31_io_in_inv_sum),
    .io_in_stage(local_pes_13_31_io_in_stage),
    .io_out_q(local_pes_13_31_io_out_q),
    .io_out_sum(local_pes_13_31_io_out_sum),
    .io_out_sum_exp(local_pes_13_31_io_out_sum_exp),
    .io_out_kv(local_pes_13_31_io_out_kv),
    .io_out_stage(local_pes_13_31_io_out_stage)
  );
  PE local_pes_14_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_0_clock),
    .reset(local_pes_14_0_reset),
    .io_in_q(local_pes_14_0_io_in_q),
    .io_in_kv(local_pes_14_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_0_io_in_inv_sum),
    .io_in_stage(local_pes_14_0_io_in_stage),
    .io_out_q(local_pes_14_0_io_out_q),
    .io_out_sum(local_pes_14_0_io_out_sum),
    .io_out_kv(local_pes_14_0_io_out_kv),
    .io_out_stage(local_pes_14_0_io_out_stage)
  );
  PE_1 local_pes_14_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_1_clock),
    .reset(local_pes_14_1_reset),
    .io_in_q(local_pes_14_1_io_in_q),
    .io_in_sum(local_pes_14_1_io_in_sum),
    .io_in_sum_exp(local_pes_14_1_io_in_sum_exp),
    .io_in_kv(local_pes_14_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_1_io_in_inv_sum),
    .io_in_stage(local_pes_14_1_io_in_stage),
    .io_out_q(local_pes_14_1_io_out_q),
    .io_out_sum(local_pes_14_1_io_out_sum),
    .io_out_sum_exp(local_pes_14_1_io_out_sum_exp),
    .io_out_kv(local_pes_14_1_io_out_kv),
    .io_out_stage(local_pes_14_1_io_out_stage)
  );
  PE_1 local_pes_14_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_2_clock),
    .reset(local_pes_14_2_reset),
    .io_in_q(local_pes_14_2_io_in_q),
    .io_in_sum(local_pes_14_2_io_in_sum),
    .io_in_sum_exp(local_pes_14_2_io_in_sum_exp),
    .io_in_kv(local_pes_14_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_2_io_in_inv_sum),
    .io_in_stage(local_pes_14_2_io_in_stage),
    .io_out_q(local_pes_14_2_io_out_q),
    .io_out_sum(local_pes_14_2_io_out_sum),
    .io_out_sum_exp(local_pes_14_2_io_out_sum_exp),
    .io_out_kv(local_pes_14_2_io_out_kv),
    .io_out_stage(local_pes_14_2_io_out_stage)
  );
  PE_1 local_pes_14_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_3_clock),
    .reset(local_pes_14_3_reset),
    .io_in_q(local_pes_14_3_io_in_q),
    .io_in_sum(local_pes_14_3_io_in_sum),
    .io_in_sum_exp(local_pes_14_3_io_in_sum_exp),
    .io_in_kv(local_pes_14_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_3_io_in_inv_sum),
    .io_in_stage(local_pes_14_3_io_in_stage),
    .io_out_q(local_pes_14_3_io_out_q),
    .io_out_sum(local_pes_14_3_io_out_sum),
    .io_out_sum_exp(local_pes_14_3_io_out_sum_exp),
    .io_out_kv(local_pes_14_3_io_out_kv),
    .io_out_stage(local_pes_14_3_io_out_stage)
  );
  PE_1 local_pes_14_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_4_clock),
    .reset(local_pes_14_4_reset),
    .io_in_q(local_pes_14_4_io_in_q),
    .io_in_sum(local_pes_14_4_io_in_sum),
    .io_in_sum_exp(local_pes_14_4_io_in_sum_exp),
    .io_in_kv(local_pes_14_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_4_io_in_inv_sum),
    .io_in_stage(local_pes_14_4_io_in_stage),
    .io_out_q(local_pes_14_4_io_out_q),
    .io_out_sum(local_pes_14_4_io_out_sum),
    .io_out_sum_exp(local_pes_14_4_io_out_sum_exp),
    .io_out_kv(local_pes_14_4_io_out_kv),
    .io_out_stage(local_pes_14_4_io_out_stage)
  );
  PE_1 local_pes_14_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_5_clock),
    .reset(local_pes_14_5_reset),
    .io_in_q(local_pes_14_5_io_in_q),
    .io_in_sum(local_pes_14_5_io_in_sum),
    .io_in_sum_exp(local_pes_14_5_io_in_sum_exp),
    .io_in_kv(local_pes_14_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_5_io_in_inv_sum),
    .io_in_stage(local_pes_14_5_io_in_stage),
    .io_out_q(local_pes_14_5_io_out_q),
    .io_out_sum(local_pes_14_5_io_out_sum),
    .io_out_sum_exp(local_pes_14_5_io_out_sum_exp),
    .io_out_kv(local_pes_14_5_io_out_kv),
    .io_out_stage(local_pes_14_5_io_out_stage)
  );
  PE_1 local_pes_14_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_6_clock),
    .reset(local_pes_14_6_reset),
    .io_in_q(local_pes_14_6_io_in_q),
    .io_in_sum(local_pes_14_6_io_in_sum),
    .io_in_sum_exp(local_pes_14_6_io_in_sum_exp),
    .io_in_kv(local_pes_14_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_6_io_in_inv_sum),
    .io_in_stage(local_pes_14_6_io_in_stage),
    .io_out_q(local_pes_14_6_io_out_q),
    .io_out_sum(local_pes_14_6_io_out_sum),
    .io_out_sum_exp(local_pes_14_6_io_out_sum_exp),
    .io_out_kv(local_pes_14_6_io_out_kv),
    .io_out_stage(local_pes_14_6_io_out_stage)
  );
  PE_1 local_pes_14_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_7_clock),
    .reset(local_pes_14_7_reset),
    .io_in_q(local_pes_14_7_io_in_q),
    .io_in_sum(local_pes_14_7_io_in_sum),
    .io_in_sum_exp(local_pes_14_7_io_in_sum_exp),
    .io_in_kv(local_pes_14_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_7_io_in_inv_sum),
    .io_in_stage(local_pes_14_7_io_in_stage),
    .io_out_q(local_pes_14_7_io_out_q),
    .io_out_sum(local_pes_14_7_io_out_sum),
    .io_out_sum_exp(local_pes_14_7_io_out_sum_exp),
    .io_out_kv(local_pes_14_7_io_out_kv),
    .io_out_stage(local_pes_14_7_io_out_stage)
  );
  PE_1 local_pes_14_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_8_clock),
    .reset(local_pes_14_8_reset),
    .io_in_q(local_pes_14_8_io_in_q),
    .io_in_sum(local_pes_14_8_io_in_sum),
    .io_in_sum_exp(local_pes_14_8_io_in_sum_exp),
    .io_in_kv(local_pes_14_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_8_io_in_inv_sum),
    .io_in_stage(local_pes_14_8_io_in_stage),
    .io_out_q(local_pes_14_8_io_out_q),
    .io_out_sum(local_pes_14_8_io_out_sum),
    .io_out_sum_exp(local_pes_14_8_io_out_sum_exp),
    .io_out_kv(local_pes_14_8_io_out_kv),
    .io_out_stage(local_pes_14_8_io_out_stage)
  );
  PE_1 local_pes_14_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_9_clock),
    .reset(local_pes_14_9_reset),
    .io_in_q(local_pes_14_9_io_in_q),
    .io_in_sum(local_pes_14_9_io_in_sum),
    .io_in_sum_exp(local_pes_14_9_io_in_sum_exp),
    .io_in_kv(local_pes_14_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_9_io_in_inv_sum),
    .io_in_stage(local_pes_14_9_io_in_stage),
    .io_out_q(local_pes_14_9_io_out_q),
    .io_out_sum(local_pes_14_9_io_out_sum),
    .io_out_sum_exp(local_pes_14_9_io_out_sum_exp),
    .io_out_kv(local_pes_14_9_io_out_kv),
    .io_out_stage(local_pes_14_9_io_out_stage)
  );
  PE_1 local_pes_14_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_10_clock),
    .reset(local_pes_14_10_reset),
    .io_in_q(local_pes_14_10_io_in_q),
    .io_in_sum(local_pes_14_10_io_in_sum),
    .io_in_sum_exp(local_pes_14_10_io_in_sum_exp),
    .io_in_kv(local_pes_14_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_10_io_in_inv_sum),
    .io_in_stage(local_pes_14_10_io_in_stage),
    .io_out_q(local_pes_14_10_io_out_q),
    .io_out_sum(local_pes_14_10_io_out_sum),
    .io_out_sum_exp(local_pes_14_10_io_out_sum_exp),
    .io_out_kv(local_pes_14_10_io_out_kv),
    .io_out_stage(local_pes_14_10_io_out_stage)
  );
  PE_1 local_pes_14_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_11_clock),
    .reset(local_pes_14_11_reset),
    .io_in_q(local_pes_14_11_io_in_q),
    .io_in_sum(local_pes_14_11_io_in_sum),
    .io_in_sum_exp(local_pes_14_11_io_in_sum_exp),
    .io_in_kv(local_pes_14_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_11_io_in_inv_sum),
    .io_in_stage(local_pes_14_11_io_in_stage),
    .io_out_q(local_pes_14_11_io_out_q),
    .io_out_sum(local_pes_14_11_io_out_sum),
    .io_out_sum_exp(local_pes_14_11_io_out_sum_exp),
    .io_out_kv(local_pes_14_11_io_out_kv),
    .io_out_stage(local_pes_14_11_io_out_stage)
  );
  PE_1 local_pes_14_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_12_clock),
    .reset(local_pes_14_12_reset),
    .io_in_q(local_pes_14_12_io_in_q),
    .io_in_sum(local_pes_14_12_io_in_sum),
    .io_in_sum_exp(local_pes_14_12_io_in_sum_exp),
    .io_in_kv(local_pes_14_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_12_io_in_inv_sum),
    .io_in_stage(local_pes_14_12_io_in_stage),
    .io_out_q(local_pes_14_12_io_out_q),
    .io_out_sum(local_pes_14_12_io_out_sum),
    .io_out_sum_exp(local_pes_14_12_io_out_sum_exp),
    .io_out_kv(local_pes_14_12_io_out_kv),
    .io_out_stage(local_pes_14_12_io_out_stage)
  );
  PE_1 local_pes_14_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_13_clock),
    .reset(local_pes_14_13_reset),
    .io_in_q(local_pes_14_13_io_in_q),
    .io_in_sum(local_pes_14_13_io_in_sum),
    .io_in_sum_exp(local_pes_14_13_io_in_sum_exp),
    .io_in_kv(local_pes_14_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_13_io_in_inv_sum),
    .io_in_stage(local_pes_14_13_io_in_stage),
    .io_out_q(local_pes_14_13_io_out_q),
    .io_out_sum(local_pes_14_13_io_out_sum),
    .io_out_sum_exp(local_pes_14_13_io_out_sum_exp),
    .io_out_kv(local_pes_14_13_io_out_kv),
    .io_out_stage(local_pes_14_13_io_out_stage)
  );
  PE_1 local_pes_14_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_14_clock),
    .reset(local_pes_14_14_reset),
    .io_in_q(local_pes_14_14_io_in_q),
    .io_in_sum(local_pes_14_14_io_in_sum),
    .io_in_sum_exp(local_pes_14_14_io_in_sum_exp),
    .io_in_kv(local_pes_14_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_14_io_in_inv_sum),
    .io_in_stage(local_pes_14_14_io_in_stage),
    .io_out_q(local_pes_14_14_io_out_q),
    .io_out_sum(local_pes_14_14_io_out_sum),
    .io_out_sum_exp(local_pes_14_14_io_out_sum_exp),
    .io_out_kv(local_pes_14_14_io_out_kv),
    .io_out_stage(local_pes_14_14_io_out_stage)
  );
  PE_1 local_pes_14_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_15_clock),
    .reset(local_pes_14_15_reset),
    .io_in_q(local_pes_14_15_io_in_q),
    .io_in_sum(local_pes_14_15_io_in_sum),
    .io_in_sum_exp(local_pes_14_15_io_in_sum_exp),
    .io_in_kv(local_pes_14_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_15_io_in_inv_sum),
    .io_in_stage(local_pes_14_15_io_in_stage),
    .io_out_q(local_pes_14_15_io_out_q),
    .io_out_sum(local_pes_14_15_io_out_sum),
    .io_out_sum_exp(local_pes_14_15_io_out_sum_exp),
    .io_out_kv(local_pes_14_15_io_out_kv),
    .io_out_stage(local_pes_14_15_io_out_stage)
  );
  PE_1 local_pes_14_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_16_clock),
    .reset(local_pes_14_16_reset),
    .io_in_q(local_pes_14_16_io_in_q),
    .io_in_sum(local_pes_14_16_io_in_sum),
    .io_in_sum_exp(local_pes_14_16_io_in_sum_exp),
    .io_in_kv(local_pes_14_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_16_io_in_inv_sum),
    .io_in_stage(local_pes_14_16_io_in_stage),
    .io_out_q(local_pes_14_16_io_out_q),
    .io_out_sum(local_pes_14_16_io_out_sum),
    .io_out_sum_exp(local_pes_14_16_io_out_sum_exp),
    .io_out_kv(local_pes_14_16_io_out_kv),
    .io_out_stage(local_pes_14_16_io_out_stage)
  );
  PE_1 local_pes_14_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_17_clock),
    .reset(local_pes_14_17_reset),
    .io_in_q(local_pes_14_17_io_in_q),
    .io_in_sum(local_pes_14_17_io_in_sum),
    .io_in_sum_exp(local_pes_14_17_io_in_sum_exp),
    .io_in_kv(local_pes_14_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_17_io_in_inv_sum),
    .io_in_stage(local_pes_14_17_io_in_stage),
    .io_out_q(local_pes_14_17_io_out_q),
    .io_out_sum(local_pes_14_17_io_out_sum),
    .io_out_sum_exp(local_pes_14_17_io_out_sum_exp),
    .io_out_kv(local_pes_14_17_io_out_kv),
    .io_out_stage(local_pes_14_17_io_out_stage)
  );
  PE_1 local_pes_14_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_18_clock),
    .reset(local_pes_14_18_reset),
    .io_in_q(local_pes_14_18_io_in_q),
    .io_in_sum(local_pes_14_18_io_in_sum),
    .io_in_sum_exp(local_pes_14_18_io_in_sum_exp),
    .io_in_kv(local_pes_14_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_18_io_in_inv_sum),
    .io_in_stage(local_pes_14_18_io_in_stage),
    .io_out_q(local_pes_14_18_io_out_q),
    .io_out_sum(local_pes_14_18_io_out_sum),
    .io_out_sum_exp(local_pes_14_18_io_out_sum_exp),
    .io_out_kv(local_pes_14_18_io_out_kv),
    .io_out_stage(local_pes_14_18_io_out_stage)
  );
  PE_1 local_pes_14_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_19_clock),
    .reset(local_pes_14_19_reset),
    .io_in_q(local_pes_14_19_io_in_q),
    .io_in_sum(local_pes_14_19_io_in_sum),
    .io_in_sum_exp(local_pes_14_19_io_in_sum_exp),
    .io_in_kv(local_pes_14_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_19_io_in_inv_sum),
    .io_in_stage(local_pes_14_19_io_in_stage),
    .io_out_q(local_pes_14_19_io_out_q),
    .io_out_sum(local_pes_14_19_io_out_sum),
    .io_out_sum_exp(local_pes_14_19_io_out_sum_exp),
    .io_out_kv(local_pes_14_19_io_out_kv),
    .io_out_stage(local_pes_14_19_io_out_stage)
  );
  PE_1 local_pes_14_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_20_clock),
    .reset(local_pes_14_20_reset),
    .io_in_q(local_pes_14_20_io_in_q),
    .io_in_sum(local_pes_14_20_io_in_sum),
    .io_in_sum_exp(local_pes_14_20_io_in_sum_exp),
    .io_in_kv(local_pes_14_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_20_io_in_inv_sum),
    .io_in_stage(local_pes_14_20_io_in_stage),
    .io_out_q(local_pes_14_20_io_out_q),
    .io_out_sum(local_pes_14_20_io_out_sum),
    .io_out_sum_exp(local_pes_14_20_io_out_sum_exp),
    .io_out_kv(local_pes_14_20_io_out_kv),
    .io_out_stage(local_pes_14_20_io_out_stage)
  );
  PE_1 local_pes_14_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_21_clock),
    .reset(local_pes_14_21_reset),
    .io_in_q(local_pes_14_21_io_in_q),
    .io_in_sum(local_pes_14_21_io_in_sum),
    .io_in_sum_exp(local_pes_14_21_io_in_sum_exp),
    .io_in_kv(local_pes_14_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_21_io_in_inv_sum),
    .io_in_stage(local_pes_14_21_io_in_stage),
    .io_out_q(local_pes_14_21_io_out_q),
    .io_out_sum(local_pes_14_21_io_out_sum),
    .io_out_sum_exp(local_pes_14_21_io_out_sum_exp),
    .io_out_kv(local_pes_14_21_io_out_kv),
    .io_out_stage(local_pes_14_21_io_out_stage)
  );
  PE_1 local_pes_14_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_22_clock),
    .reset(local_pes_14_22_reset),
    .io_in_q(local_pes_14_22_io_in_q),
    .io_in_sum(local_pes_14_22_io_in_sum),
    .io_in_sum_exp(local_pes_14_22_io_in_sum_exp),
    .io_in_kv(local_pes_14_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_22_io_in_inv_sum),
    .io_in_stage(local_pes_14_22_io_in_stage),
    .io_out_q(local_pes_14_22_io_out_q),
    .io_out_sum(local_pes_14_22_io_out_sum),
    .io_out_sum_exp(local_pes_14_22_io_out_sum_exp),
    .io_out_kv(local_pes_14_22_io_out_kv),
    .io_out_stage(local_pes_14_22_io_out_stage)
  );
  PE_1 local_pes_14_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_23_clock),
    .reset(local_pes_14_23_reset),
    .io_in_q(local_pes_14_23_io_in_q),
    .io_in_sum(local_pes_14_23_io_in_sum),
    .io_in_sum_exp(local_pes_14_23_io_in_sum_exp),
    .io_in_kv(local_pes_14_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_23_io_in_inv_sum),
    .io_in_stage(local_pes_14_23_io_in_stage),
    .io_out_q(local_pes_14_23_io_out_q),
    .io_out_sum(local_pes_14_23_io_out_sum),
    .io_out_sum_exp(local_pes_14_23_io_out_sum_exp),
    .io_out_kv(local_pes_14_23_io_out_kv),
    .io_out_stage(local_pes_14_23_io_out_stage)
  );
  PE_1 local_pes_14_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_24_clock),
    .reset(local_pes_14_24_reset),
    .io_in_q(local_pes_14_24_io_in_q),
    .io_in_sum(local_pes_14_24_io_in_sum),
    .io_in_sum_exp(local_pes_14_24_io_in_sum_exp),
    .io_in_kv(local_pes_14_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_24_io_in_inv_sum),
    .io_in_stage(local_pes_14_24_io_in_stage),
    .io_out_q(local_pes_14_24_io_out_q),
    .io_out_sum(local_pes_14_24_io_out_sum),
    .io_out_sum_exp(local_pes_14_24_io_out_sum_exp),
    .io_out_kv(local_pes_14_24_io_out_kv),
    .io_out_stage(local_pes_14_24_io_out_stage)
  );
  PE_1 local_pes_14_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_25_clock),
    .reset(local_pes_14_25_reset),
    .io_in_q(local_pes_14_25_io_in_q),
    .io_in_sum(local_pes_14_25_io_in_sum),
    .io_in_sum_exp(local_pes_14_25_io_in_sum_exp),
    .io_in_kv(local_pes_14_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_25_io_in_inv_sum),
    .io_in_stage(local_pes_14_25_io_in_stage),
    .io_out_q(local_pes_14_25_io_out_q),
    .io_out_sum(local_pes_14_25_io_out_sum),
    .io_out_sum_exp(local_pes_14_25_io_out_sum_exp),
    .io_out_kv(local_pes_14_25_io_out_kv),
    .io_out_stage(local_pes_14_25_io_out_stage)
  );
  PE_1 local_pes_14_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_26_clock),
    .reset(local_pes_14_26_reset),
    .io_in_q(local_pes_14_26_io_in_q),
    .io_in_sum(local_pes_14_26_io_in_sum),
    .io_in_sum_exp(local_pes_14_26_io_in_sum_exp),
    .io_in_kv(local_pes_14_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_26_io_in_inv_sum),
    .io_in_stage(local_pes_14_26_io_in_stage),
    .io_out_q(local_pes_14_26_io_out_q),
    .io_out_sum(local_pes_14_26_io_out_sum),
    .io_out_sum_exp(local_pes_14_26_io_out_sum_exp),
    .io_out_kv(local_pes_14_26_io_out_kv),
    .io_out_stage(local_pes_14_26_io_out_stage)
  );
  PE_1 local_pes_14_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_27_clock),
    .reset(local_pes_14_27_reset),
    .io_in_q(local_pes_14_27_io_in_q),
    .io_in_sum(local_pes_14_27_io_in_sum),
    .io_in_sum_exp(local_pes_14_27_io_in_sum_exp),
    .io_in_kv(local_pes_14_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_27_io_in_inv_sum),
    .io_in_stage(local_pes_14_27_io_in_stage),
    .io_out_q(local_pes_14_27_io_out_q),
    .io_out_sum(local_pes_14_27_io_out_sum),
    .io_out_sum_exp(local_pes_14_27_io_out_sum_exp),
    .io_out_kv(local_pes_14_27_io_out_kv),
    .io_out_stage(local_pes_14_27_io_out_stage)
  );
  PE_1 local_pes_14_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_28_clock),
    .reset(local_pes_14_28_reset),
    .io_in_q(local_pes_14_28_io_in_q),
    .io_in_sum(local_pes_14_28_io_in_sum),
    .io_in_sum_exp(local_pes_14_28_io_in_sum_exp),
    .io_in_kv(local_pes_14_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_28_io_in_inv_sum),
    .io_in_stage(local_pes_14_28_io_in_stage),
    .io_out_q(local_pes_14_28_io_out_q),
    .io_out_sum(local_pes_14_28_io_out_sum),
    .io_out_sum_exp(local_pes_14_28_io_out_sum_exp),
    .io_out_kv(local_pes_14_28_io_out_kv),
    .io_out_stage(local_pes_14_28_io_out_stage)
  );
  PE_1 local_pes_14_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_29_clock),
    .reset(local_pes_14_29_reset),
    .io_in_q(local_pes_14_29_io_in_q),
    .io_in_sum(local_pes_14_29_io_in_sum),
    .io_in_sum_exp(local_pes_14_29_io_in_sum_exp),
    .io_in_kv(local_pes_14_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_29_io_in_inv_sum),
    .io_in_stage(local_pes_14_29_io_in_stage),
    .io_out_q(local_pes_14_29_io_out_q),
    .io_out_sum(local_pes_14_29_io_out_sum),
    .io_out_sum_exp(local_pes_14_29_io_out_sum_exp),
    .io_out_kv(local_pes_14_29_io_out_kv),
    .io_out_stage(local_pes_14_29_io_out_stage)
  );
  PE_1 local_pes_14_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_30_clock),
    .reset(local_pes_14_30_reset),
    .io_in_q(local_pes_14_30_io_in_q),
    .io_in_sum(local_pes_14_30_io_in_sum),
    .io_in_sum_exp(local_pes_14_30_io_in_sum_exp),
    .io_in_kv(local_pes_14_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_30_io_in_inv_sum),
    .io_in_stage(local_pes_14_30_io_in_stage),
    .io_out_q(local_pes_14_30_io_out_q),
    .io_out_sum(local_pes_14_30_io_out_sum),
    .io_out_sum_exp(local_pes_14_30_io_out_sum_exp),
    .io_out_kv(local_pes_14_30_io_out_kv),
    .io_out_stage(local_pes_14_30_io_out_stage)
  );
  PE_1 local_pes_14_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_14_31_clock),
    .reset(local_pes_14_31_reset),
    .io_in_q(local_pes_14_31_io_in_q),
    .io_in_sum(local_pes_14_31_io_in_sum),
    .io_in_sum_exp(local_pes_14_31_io_in_sum_exp),
    .io_in_kv(local_pes_14_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_14_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_14_31_io_in_inv_sum),
    .io_in_stage(local_pes_14_31_io_in_stage),
    .io_out_q(local_pes_14_31_io_out_q),
    .io_out_sum(local_pes_14_31_io_out_sum),
    .io_out_sum_exp(local_pes_14_31_io_out_sum_exp),
    .io_out_kv(local_pes_14_31_io_out_kv),
    .io_out_stage(local_pes_14_31_io_out_stage)
  );
  PE local_pes_15_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_0_clock),
    .reset(local_pes_15_0_reset),
    .io_in_q(local_pes_15_0_io_in_q),
    .io_in_kv(local_pes_15_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_0_io_in_inv_sum),
    .io_in_stage(local_pes_15_0_io_in_stage),
    .io_out_q(local_pes_15_0_io_out_q),
    .io_out_sum(local_pes_15_0_io_out_sum),
    .io_out_kv(local_pes_15_0_io_out_kv),
    .io_out_stage(local_pes_15_0_io_out_stage)
  );
  PE_1 local_pes_15_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_1_clock),
    .reset(local_pes_15_1_reset),
    .io_in_q(local_pes_15_1_io_in_q),
    .io_in_sum(local_pes_15_1_io_in_sum),
    .io_in_sum_exp(local_pes_15_1_io_in_sum_exp),
    .io_in_kv(local_pes_15_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_1_io_in_inv_sum),
    .io_in_stage(local_pes_15_1_io_in_stage),
    .io_out_q(local_pes_15_1_io_out_q),
    .io_out_sum(local_pes_15_1_io_out_sum),
    .io_out_sum_exp(local_pes_15_1_io_out_sum_exp),
    .io_out_kv(local_pes_15_1_io_out_kv),
    .io_out_stage(local_pes_15_1_io_out_stage)
  );
  PE_1 local_pes_15_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_2_clock),
    .reset(local_pes_15_2_reset),
    .io_in_q(local_pes_15_2_io_in_q),
    .io_in_sum(local_pes_15_2_io_in_sum),
    .io_in_sum_exp(local_pes_15_2_io_in_sum_exp),
    .io_in_kv(local_pes_15_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_2_io_in_inv_sum),
    .io_in_stage(local_pes_15_2_io_in_stage),
    .io_out_q(local_pes_15_2_io_out_q),
    .io_out_sum(local_pes_15_2_io_out_sum),
    .io_out_sum_exp(local_pes_15_2_io_out_sum_exp),
    .io_out_kv(local_pes_15_2_io_out_kv),
    .io_out_stage(local_pes_15_2_io_out_stage)
  );
  PE_1 local_pes_15_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_3_clock),
    .reset(local_pes_15_3_reset),
    .io_in_q(local_pes_15_3_io_in_q),
    .io_in_sum(local_pes_15_3_io_in_sum),
    .io_in_sum_exp(local_pes_15_3_io_in_sum_exp),
    .io_in_kv(local_pes_15_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_3_io_in_inv_sum),
    .io_in_stage(local_pes_15_3_io_in_stage),
    .io_out_q(local_pes_15_3_io_out_q),
    .io_out_sum(local_pes_15_3_io_out_sum),
    .io_out_sum_exp(local_pes_15_3_io_out_sum_exp),
    .io_out_kv(local_pes_15_3_io_out_kv),
    .io_out_stage(local_pes_15_3_io_out_stage)
  );
  PE_1 local_pes_15_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_4_clock),
    .reset(local_pes_15_4_reset),
    .io_in_q(local_pes_15_4_io_in_q),
    .io_in_sum(local_pes_15_4_io_in_sum),
    .io_in_sum_exp(local_pes_15_4_io_in_sum_exp),
    .io_in_kv(local_pes_15_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_4_io_in_inv_sum),
    .io_in_stage(local_pes_15_4_io_in_stage),
    .io_out_q(local_pes_15_4_io_out_q),
    .io_out_sum(local_pes_15_4_io_out_sum),
    .io_out_sum_exp(local_pes_15_4_io_out_sum_exp),
    .io_out_kv(local_pes_15_4_io_out_kv),
    .io_out_stage(local_pes_15_4_io_out_stage)
  );
  PE_1 local_pes_15_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_5_clock),
    .reset(local_pes_15_5_reset),
    .io_in_q(local_pes_15_5_io_in_q),
    .io_in_sum(local_pes_15_5_io_in_sum),
    .io_in_sum_exp(local_pes_15_5_io_in_sum_exp),
    .io_in_kv(local_pes_15_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_5_io_in_inv_sum),
    .io_in_stage(local_pes_15_5_io_in_stage),
    .io_out_q(local_pes_15_5_io_out_q),
    .io_out_sum(local_pes_15_5_io_out_sum),
    .io_out_sum_exp(local_pes_15_5_io_out_sum_exp),
    .io_out_kv(local_pes_15_5_io_out_kv),
    .io_out_stage(local_pes_15_5_io_out_stage)
  );
  PE_1 local_pes_15_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_6_clock),
    .reset(local_pes_15_6_reset),
    .io_in_q(local_pes_15_6_io_in_q),
    .io_in_sum(local_pes_15_6_io_in_sum),
    .io_in_sum_exp(local_pes_15_6_io_in_sum_exp),
    .io_in_kv(local_pes_15_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_6_io_in_inv_sum),
    .io_in_stage(local_pes_15_6_io_in_stage),
    .io_out_q(local_pes_15_6_io_out_q),
    .io_out_sum(local_pes_15_6_io_out_sum),
    .io_out_sum_exp(local_pes_15_6_io_out_sum_exp),
    .io_out_kv(local_pes_15_6_io_out_kv),
    .io_out_stage(local_pes_15_6_io_out_stage)
  );
  PE_1 local_pes_15_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_7_clock),
    .reset(local_pes_15_7_reset),
    .io_in_q(local_pes_15_7_io_in_q),
    .io_in_sum(local_pes_15_7_io_in_sum),
    .io_in_sum_exp(local_pes_15_7_io_in_sum_exp),
    .io_in_kv(local_pes_15_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_7_io_in_inv_sum),
    .io_in_stage(local_pes_15_7_io_in_stage),
    .io_out_q(local_pes_15_7_io_out_q),
    .io_out_sum(local_pes_15_7_io_out_sum),
    .io_out_sum_exp(local_pes_15_7_io_out_sum_exp),
    .io_out_kv(local_pes_15_7_io_out_kv),
    .io_out_stage(local_pes_15_7_io_out_stage)
  );
  PE_1 local_pes_15_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_8_clock),
    .reset(local_pes_15_8_reset),
    .io_in_q(local_pes_15_8_io_in_q),
    .io_in_sum(local_pes_15_8_io_in_sum),
    .io_in_sum_exp(local_pes_15_8_io_in_sum_exp),
    .io_in_kv(local_pes_15_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_8_io_in_inv_sum),
    .io_in_stage(local_pes_15_8_io_in_stage),
    .io_out_q(local_pes_15_8_io_out_q),
    .io_out_sum(local_pes_15_8_io_out_sum),
    .io_out_sum_exp(local_pes_15_8_io_out_sum_exp),
    .io_out_kv(local_pes_15_8_io_out_kv),
    .io_out_stage(local_pes_15_8_io_out_stage)
  );
  PE_1 local_pes_15_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_9_clock),
    .reset(local_pes_15_9_reset),
    .io_in_q(local_pes_15_9_io_in_q),
    .io_in_sum(local_pes_15_9_io_in_sum),
    .io_in_sum_exp(local_pes_15_9_io_in_sum_exp),
    .io_in_kv(local_pes_15_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_9_io_in_inv_sum),
    .io_in_stage(local_pes_15_9_io_in_stage),
    .io_out_q(local_pes_15_9_io_out_q),
    .io_out_sum(local_pes_15_9_io_out_sum),
    .io_out_sum_exp(local_pes_15_9_io_out_sum_exp),
    .io_out_kv(local_pes_15_9_io_out_kv),
    .io_out_stage(local_pes_15_9_io_out_stage)
  );
  PE_1 local_pes_15_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_10_clock),
    .reset(local_pes_15_10_reset),
    .io_in_q(local_pes_15_10_io_in_q),
    .io_in_sum(local_pes_15_10_io_in_sum),
    .io_in_sum_exp(local_pes_15_10_io_in_sum_exp),
    .io_in_kv(local_pes_15_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_10_io_in_inv_sum),
    .io_in_stage(local_pes_15_10_io_in_stage),
    .io_out_q(local_pes_15_10_io_out_q),
    .io_out_sum(local_pes_15_10_io_out_sum),
    .io_out_sum_exp(local_pes_15_10_io_out_sum_exp),
    .io_out_kv(local_pes_15_10_io_out_kv),
    .io_out_stage(local_pes_15_10_io_out_stage)
  );
  PE_1 local_pes_15_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_11_clock),
    .reset(local_pes_15_11_reset),
    .io_in_q(local_pes_15_11_io_in_q),
    .io_in_sum(local_pes_15_11_io_in_sum),
    .io_in_sum_exp(local_pes_15_11_io_in_sum_exp),
    .io_in_kv(local_pes_15_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_11_io_in_inv_sum),
    .io_in_stage(local_pes_15_11_io_in_stage),
    .io_out_q(local_pes_15_11_io_out_q),
    .io_out_sum(local_pes_15_11_io_out_sum),
    .io_out_sum_exp(local_pes_15_11_io_out_sum_exp),
    .io_out_kv(local_pes_15_11_io_out_kv),
    .io_out_stage(local_pes_15_11_io_out_stage)
  );
  PE_1 local_pes_15_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_12_clock),
    .reset(local_pes_15_12_reset),
    .io_in_q(local_pes_15_12_io_in_q),
    .io_in_sum(local_pes_15_12_io_in_sum),
    .io_in_sum_exp(local_pes_15_12_io_in_sum_exp),
    .io_in_kv(local_pes_15_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_12_io_in_inv_sum),
    .io_in_stage(local_pes_15_12_io_in_stage),
    .io_out_q(local_pes_15_12_io_out_q),
    .io_out_sum(local_pes_15_12_io_out_sum),
    .io_out_sum_exp(local_pes_15_12_io_out_sum_exp),
    .io_out_kv(local_pes_15_12_io_out_kv),
    .io_out_stage(local_pes_15_12_io_out_stage)
  );
  PE_1 local_pes_15_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_13_clock),
    .reset(local_pes_15_13_reset),
    .io_in_q(local_pes_15_13_io_in_q),
    .io_in_sum(local_pes_15_13_io_in_sum),
    .io_in_sum_exp(local_pes_15_13_io_in_sum_exp),
    .io_in_kv(local_pes_15_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_13_io_in_inv_sum),
    .io_in_stage(local_pes_15_13_io_in_stage),
    .io_out_q(local_pes_15_13_io_out_q),
    .io_out_sum(local_pes_15_13_io_out_sum),
    .io_out_sum_exp(local_pes_15_13_io_out_sum_exp),
    .io_out_kv(local_pes_15_13_io_out_kv),
    .io_out_stage(local_pes_15_13_io_out_stage)
  );
  PE_1 local_pes_15_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_14_clock),
    .reset(local_pes_15_14_reset),
    .io_in_q(local_pes_15_14_io_in_q),
    .io_in_sum(local_pes_15_14_io_in_sum),
    .io_in_sum_exp(local_pes_15_14_io_in_sum_exp),
    .io_in_kv(local_pes_15_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_14_io_in_inv_sum),
    .io_in_stage(local_pes_15_14_io_in_stage),
    .io_out_q(local_pes_15_14_io_out_q),
    .io_out_sum(local_pes_15_14_io_out_sum),
    .io_out_sum_exp(local_pes_15_14_io_out_sum_exp),
    .io_out_kv(local_pes_15_14_io_out_kv),
    .io_out_stage(local_pes_15_14_io_out_stage)
  );
  PE_1 local_pes_15_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_15_clock),
    .reset(local_pes_15_15_reset),
    .io_in_q(local_pes_15_15_io_in_q),
    .io_in_sum(local_pes_15_15_io_in_sum),
    .io_in_sum_exp(local_pes_15_15_io_in_sum_exp),
    .io_in_kv(local_pes_15_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_15_io_in_inv_sum),
    .io_in_stage(local_pes_15_15_io_in_stage),
    .io_out_q(local_pes_15_15_io_out_q),
    .io_out_sum(local_pes_15_15_io_out_sum),
    .io_out_sum_exp(local_pes_15_15_io_out_sum_exp),
    .io_out_kv(local_pes_15_15_io_out_kv),
    .io_out_stage(local_pes_15_15_io_out_stage)
  );
  PE_1 local_pes_15_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_16_clock),
    .reset(local_pes_15_16_reset),
    .io_in_q(local_pes_15_16_io_in_q),
    .io_in_sum(local_pes_15_16_io_in_sum),
    .io_in_sum_exp(local_pes_15_16_io_in_sum_exp),
    .io_in_kv(local_pes_15_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_16_io_in_inv_sum),
    .io_in_stage(local_pes_15_16_io_in_stage),
    .io_out_q(local_pes_15_16_io_out_q),
    .io_out_sum(local_pes_15_16_io_out_sum),
    .io_out_sum_exp(local_pes_15_16_io_out_sum_exp),
    .io_out_kv(local_pes_15_16_io_out_kv),
    .io_out_stage(local_pes_15_16_io_out_stage)
  );
  PE_1 local_pes_15_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_17_clock),
    .reset(local_pes_15_17_reset),
    .io_in_q(local_pes_15_17_io_in_q),
    .io_in_sum(local_pes_15_17_io_in_sum),
    .io_in_sum_exp(local_pes_15_17_io_in_sum_exp),
    .io_in_kv(local_pes_15_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_17_io_in_inv_sum),
    .io_in_stage(local_pes_15_17_io_in_stage),
    .io_out_q(local_pes_15_17_io_out_q),
    .io_out_sum(local_pes_15_17_io_out_sum),
    .io_out_sum_exp(local_pes_15_17_io_out_sum_exp),
    .io_out_kv(local_pes_15_17_io_out_kv),
    .io_out_stage(local_pes_15_17_io_out_stage)
  );
  PE_1 local_pes_15_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_18_clock),
    .reset(local_pes_15_18_reset),
    .io_in_q(local_pes_15_18_io_in_q),
    .io_in_sum(local_pes_15_18_io_in_sum),
    .io_in_sum_exp(local_pes_15_18_io_in_sum_exp),
    .io_in_kv(local_pes_15_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_18_io_in_inv_sum),
    .io_in_stage(local_pes_15_18_io_in_stage),
    .io_out_q(local_pes_15_18_io_out_q),
    .io_out_sum(local_pes_15_18_io_out_sum),
    .io_out_sum_exp(local_pes_15_18_io_out_sum_exp),
    .io_out_kv(local_pes_15_18_io_out_kv),
    .io_out_stage(local_pes_15_18_io_out_stage)
  );
  PE_1 local_pes_15_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_19_clock),
    .reset(local_pes_15_19_reset),
    .io_in_q(local_pes_15_19_io_in_q),
    .io_in_sum(local_pes_15_19_io_in_sum),
    .io_in_sum_exp(local_pes_15_19_io_in_sum_exp),
    .io_in_kv(local_pes_15_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_19_io_in_inv_sum),
    .io_in_stage(local_pes_15_19_io_in_stage),
    .io_out_q(local_pes_15_19_io_out_q),
    .io_out_sum(local_pes_15_19_io_out_sum),
    .io_out_sum_exp(local_pes_15_19_io_out_sum_exp),
    .io_out_kv(local_pes_15_19_io_out_kv),
    .io_out_stage(local_pes_15_19_io_out_stage)
  );
  PE_1 local_pes_15_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_20_clock),
    .reset(local_pes_15_20_reset),
    .io_in_q(local_pes_15_20_io_in_q),
    .io_in_sum(local_pes_15_20_io_in_sum),
    .io_in_sum_exp(local_pes_15_20_io_in_sum_exp),
    .io_in_kv(local_pes_15_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_20_io_in_inv_sum),
    .io_in_stage(local_pes_15_20_io_in_stage),
    .io_out_q(local_pes_15_20_io_out_q),
    .io_out_sum(local_pes_15_20_io_out_sum),
    .io_out_sum_exp(local_pes_15_20_io_out_sum_exp),
    .io_out_kv(local_pes_15_20_io_out_kv),
    .io_out_stage(local_pes_15_20_io_out_stage)
  );
  PE_1 local_pes_15_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_21_clock),
    .reset(local_pes_15_21_reset),
    .io_in_q(local_pes_15_21_io_in_q),
    .io_in_sum(local_pes_15_21_io_in_sum),
    .io_in_sum_exp(local_pes_15_21_io_in_sum_exp),
    .io_in_kv(local_pes_15_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_21_io_in_inv_sum),
    .io_in_stage(local_pes_15_21_io_in_stage),
    .io_out_q(local_pes_15_21_io_out_q),
    .io_out_sum(local_pes_15_21_io_out_sum),
    .io_out_sum_exp(local_pes_15_21_io_out_sum_exp),
    .io_out_kv(local_pes_15_21_io_out_kv),
    .io_out_stage(local_pes_15_21_io_out_stage)
  );
  PE_1 local_pes_15_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_22_clock),
    .reset(local_pes_15_22_reset),
    .io_in_q(local_pes_15_22_io_in_q),
    .io_in_sum(local_pes_15_22_io_in_sum),
    .io_in_sum_exp(local_pes_15_22_io_in_sum_exp),
    .io_in_kv(local_pes_15_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_22_io_in_inv_sum),
    .io_in_stage(local_pes_15_22_io_in_stage),
    .io_out_q(local_pes_15_22_io_out_q),
    .io_out_sum(local_pes_15_22_io_out_sum),
    .io_out_sum_exp(local_pes_15_22_io_out_sum_exp),
    .io_out_kv(local_pes_15_22_io_out_kv),
    .io_out_stage(local_pes_15_22_io_out_stage)
  );
  PE_1 local_pes_15_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_23_clock),
    .reset(local_pes_15_23_reset),
    .io_in_q(local_pes_15_23_io_in_q),
    .io_in_sum(local_pes_15_23_io_in_sum),
    .io_in_sum_exp(local_pes_15_23_io_in_sum_exp),
    .io_in_kv(local_pes_15_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_23_io_in_inv_sum),
    .io_in_stage(local_pes_15_23_io_in_stage),
    .io_out_q(local_pes_15_23_io_out_q),
    .io_out_sum(local_pes_15_23_io_out_sum),
    .io_out_sum_exp(local_pes_15_23_io_out_sum_exp),
    .io_out_kv(local_pes_15_23_io_out_kv),
    .io_out_stage(local_pes_15_23_io_out_stage)
  );
  PE_1 local_pes_15_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_24_clock),
    .reset(local_pes_15_24_reset),
    .io_in_q(local_pes_15_24_io_in_q),
    .io_in_sum(local_pes_15_24_io_in_sum),
    .io_in_sum_exp(local_pes_15_24_io_in_sum_exp),
    .io_in_kv(local_pes_15_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_24_io_in_inv_sum),
    .io_in_stage(local_pes_15_24_io_in_stage),
    .io_out_q(local_pes_15_24_io_out_q),
    .io_out_sum(local_pes_15_24_io_out_sum),
    .io_out_sum_exp(local_pes_15_24_io_out_sum_exp),
    .io_out_kv(local_pes_15_24_io_out_kv),
    .io_out_stage(local_pes_15_24_io_out_stage)
  );
  PE_1 local_pes_15_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_25_clock),
    .reset(local_pes_15_25_reset),
    .io_in_q(local_pes_15_25_io_in_q),
    .io_in_sum(local_pes_15_25_io_in_sum),
    .io_in_sum_exp(local_pes_15_25_io_in_sum_exp),
    .io_in_kv(local_pes_15_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_25_io_in_inv_sum),
    .io_in_stage(local_pes_15_25_io_in_stage),
    .io_out_q(local_pes_15_25_io_out_q),
    .io_out_sum(local_pes_15_25_io_out_sum),
    .io_out_sum_exp(local_pes_15_25_io_out_sum_exp),
    .io_out_kv(local_pes_15_25_io_out_kv),
    .io_out_stage(local_pes_15_25_io_out_stage)
  );
  PE_1 local_pes_15_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_26_clock),
    .reset(local_pes_15_26_reset),
    .io_in_q(local_pes_15_26_io_in_q),
    .io_in_sum(local_pes_15_26_io_in_sum),
    .io_in_sum_exp(local_pes_15_26_io_in_sum_exp),
    .io_in_kv(local_pes_15_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_26_io_in_inv_sum),
    .io_in_stage(local_pes_15_26_io_in_stage),
    .io_out_q(local_pes_15_26_io_out_q),
    .io_out_sum(local_pes_15_26_io_out_sum),
    .io_out_sum_exp(local_pes_15_26_io_out_sum_exp),
    .io_out_kv(local_pes_15_26_io_out_kv),
    .io_out_stage(local_pes_15_26_io_out_stage)
  );
  PE_1 local_pes_15_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_27_clock),
    .reset(local_pes_15_27_reset),
    .io_in_q(local_pes_15_27_io_in_q),
    .io_in_sum(local_pes_15_27_io_in_sum),
    .io_in_sum_exp(local_pes_15_27_io_in_sum_exp),
    .io_in_kv(local_pes_15_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_27_io_in_inv_sum),
    .io_in_stage(local_pes_15_27_io_in_stage),
    .io_out_q(local_pes_15_27_io_out_q),
    .io_out_sum(local_pes_15_27_io_out_sum),
    .io_out_sum_exp(local_pes_15_27_io_out_sum_exp),
    .io_out_kv(local_pes_15_27_io_out_kv),
    .io_out_stage(local_pes_15_27_io_out_stage)
  );
  PE_1 local_pes_15_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_28_clock),
    .reset(local_pes_15_28_reset),
    .io_in_q(local_pes_15_28_io_in_q),
    .io_in_sum(local_pes_15_28_io_in_sum),
    .io_in_sum_exp(local_pes_15_28_io_in_sum_exp),
    .io_in_kv(local_pes_15_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_28_io_in_inv_sum),
    .io_in_stage(local_pes_15_28_io_in_stage),
    .io_out_q(local_pes_15_28_io_out_q),
    .io_out_sum(local_pes_15_28_io_out_sum),
    .io_out_sum_exp(local_pes_15_28_io_out_sum_exp),
    .io_out_kv(local_pes_15_28_io_out_kv),
    .io_out_stage(local_pes_15_28_io_out_stage)
  );
  PE_1 local_pes_15_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_29_clock),
    .reset(local_pes_15_29_reset),
    .io_in_q(local_pes_15_29_io_in_q),
    .io_in_sum(local_pes_15_29_io_in_sum),
    .io_in_sum_exp(local_pes_15_29_io_in_sum_exp),
    .io_in_kv(local_pes_15_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_29_io_in_inv_sum),
    .io_in_stage(local_pes_15_29_io_in_stage),
    .io_out_q(local_pes_15_29_io_out_q),
    .io_out_sum(local_pes_15_29_io_out_sum),
    .io_out_sum_exp(local_pes_15_29_io_out_sum_exp),
    .io_out_kv(local_pes_15_29_io_out_kv),
    .io_out_stage(local_pes_15_29_io_out_stage)
  );
  PE_1 local_pes_15_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_30_clock),
    .reset(local_pes_15_30_reset),
    .io_in_q(local_pes_15_30_io_in_q),
    .io_in_sum(local_pes_15_30_io_in_sum),
    .io_in_sum_exp(local_pes_15_30_io_in_sum_exp),
    .io_in_kv(local_pes_15_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_30_io_in_inv_sum),
    .io_in_stage(local_pes_15_30_io_in_stage),
    .io_out_q(local_pes_15_30_io_out_q),
    .io_out_sum(local_pes_15_30_io_out_sum),
    .io_out_sum_exp(local_pes_15_30_io_out_sum_exp),
    .io_out_kv(local_pes_15_30_io_out_kv),
    .io_out_stage(local_pes_15_30_io_out_stage)
  );
  PE_1 local_pes_15_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_15_31_clock),
    .reset(local_pes_15_31_reset),
    .io_in_q(local_pes_15_31_io_in_q),
    .io_in_sum(local_pes_15_31_io_in_sum),
    .io_in_sum_exp(local_pes_15_31_io_in_sum_exp),
    .io_in_kv(local_pes_15_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_15_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_15_31_io_in_inv_sum),
    .io_in_stage(local_pes_15_31_io_in_stage),
    .io_out_q(local_pes_15_31_io_out_q),
    .io_out_sum(local_pes_15_31_io_out_sum),
    .io_out_sum_exp(local_pes_15_31_io_out_sum_exp),
    .io_out_kv(local_pes_15_31_io_out_kv),
    .io_out_stage(local_pes_15_31_io_out_stage)
  );
  PE local_pes_16_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_0_clock),
    .reset(local_pes_16_0_reset),
    .io_in_q(local_pes_16_0_io_in_q),
    .io_in_kv(local_pes_16_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_0_io_in_inv_sum),
    .io_in_stage(local_pes_16_0_io_in_stage),
    .io_out_q(local_pes_16_0_io_out_q),
    .io_out_sum(local_pes_16_0_io_out_sum),
    .io_out_kv(local_pes_16_0_io_out_kv),
    .io_out_stage(local_pes_16_0_io_out_stage)
  );
  PE_1 local_pes_16_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_1_clock),
    .reset(local_pes_16_1_reset),
    .io_in_q(local_pes_16_1_io_in_q),
    .io_in_sum(local_pes_16_1_io_in_sum),
    .io_in_sum_exp(local_pes_16_1_io_in_sum_exp),
    .io_in_kv(local_pes_16_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_1_io_in_inv_sum),
    .io_in_stage(local_pes_16_1_io_in_stage),
    .io_out_q(local_pes_16_1_io_out_q),
    .io_out_sum(local_pes_16_1_io_out_sum),
    .io_out_sum_exp(local_pes_16_1_io_out_sum_exp),
    .io_out_kv(local_pes_16_1_io_out_kv),
    .io_out_stage(local_pes_16_1_io_out_stage)
  );
  PE_1 local_pes_16_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_2_clock),
    .reset(local_pes_16_2_reset),
    .io_in_q(local_pes_16_2_io_in_q),
    .io_in_sum(local_pes_16_2_io_in_sum),
    .io_in_sum_exp(local_pes_16_2_io_in_sum_exp),
    .io_in_kv(local_pes_16_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_2_io_in_inv_sum),
    .io_in_stage(local_pes_16_2_io_in_stage),
    .io_out_q(local_pes_16_2_io_out_q),
    .io_out_sum(local_pes_16_2_io_out_sum),
    .io_out_sum_exp(local_pes_16_2_io_out_sum_exp),
    .io_out_kv(local_pes_16_2_io_out_kv),
    .io_out_stage(local_pes_16_2_io_out_stage)
  );
  PE_1 local_pes_16_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_3_clock),
    .reset(local_pes_16_3_reset),
    .io_in_q(local_pes_16_3_io_in_q),
    .io_in_sum(local_pes_16_3_io_in_sum),
    .io_in_sum_exp(local_pes_16_3_io_in_sum_exp),
    .io_in_kv(local_pes_16_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_3_io_in_inv_sum),
    .io_in_stage(local_pes_16_3_io_in_stage),
    .io_out_q(local_pes_16_3_io_out_q),
    .io_out_sum(local_pes_16_3_io_out_sum),
    .io_out_sum_exp(local_pes_16_3_io_out_sum_exp),
    .io_out_kv(local_pes_16_3_io_out_kv),
    .io_out_stage(local_pes_16_3_io_out_stage)
  );
  PE_1 local_pes_16_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_4_clock),
    .reset(local_pes_16_4_reset),
    .io_in_q(local_pes_16_4_io_in_q),
    .io_in_sum(local_pes_16_4_io_in_sum),
    .io_in_sum_exp(local_pes_16_4_io_in_sum_exp),
    .io_in_kv(local_pes_16_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_4_io_in_inv_sum),
    .io_in_stage(local_pes_16_4_io_in_stage),
    .io_out_q(local_pes_16_4_io_out_q),
    .io_out_sum(local_pes_16_4_io_out_sum),
    .io_out_sum_exp(local_pes_16_4_io_out_sum_exp),
    .io_out_kv(local_pes_16_4_io_out_kv),
    .io_out_stage(local_pes_16_4_io_out_stage)
  );
  PE_1 local_pes_16_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_5_clock),
    .reset(local_pes_16_5_reset),
    .io_in_q(local_pes_16_5_io_in_q),
    .io_in_sum(local_pes_16_5_io_in_sum),
    .io_in_sum_exp(local_pes_16_5_io_in_sum_exp),
    .io_in_kv(local_pes_16_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_5_io_in_inv_sum),
    .io_in_stage(local_pes_16_5_io_in_stage),
    .io_out_q(local_pes_16_5_io_out_q),
    .io_out_sum(local_pes_16_5_io_out_sum),
    .io_out_sum_exp(local_pes_16_5_io_out_sum_exp),
    .io_out_kv(local_pes_16_5_io_out_kv),
    .io_out_stage(local_pes_16_5_io_out_stage)
  );
  PE_1 local_pes_16_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_6_clock),
    .reset(local_pes_16_6_reset),
    .io_in_q(local_pes_16_6_io_in_q),
    .io_in_sum(local_pes_16_6_io_in_sum),
    .io_in_sum_exp(local_pes_16_6_io_in_sum_exp),
    .io_in_kv(local_pes_16_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_6_io_in_inv_sum),
    .io_in_stage(local_pes_16_6_io_in_stage),
    .io_out_q(local_pes_16_6_io_out_q),
    .io_out_sum(local_pes_16_6_io_out_sum),
    .io_out_sum_exp(local_pes_16_6_io_out_sum_exp),
    .io_out_kv(local_pes_16_6_io_out_kv),
    .io_out_stage(local_pes_16_6_io_out_stage)
  );
  PE_1 local_pes_16_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_7_clock),
    .reset(local_pes_16_7_reset),
    .io_in_q(local_pes_16_7_io_in_q),
    .io_in_sum(local_pes_16_7_io_in_sum),
    .io_in_sum_exp(local_pes_16_7_io_in_sum_exp),
    .io_in_kv(local_pes_16_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_7_io_in_inv_sum),
    .io_in_stage(local_pes_16_7_io_in_stage),
    .io_out_q(local_pes_16_7_io_out_q),
    .io_out_sum(local_pes_16_7_io_out_sum),
    .io_out_sum_exp(local_pes_16_7_io_out_sum_exp),
    .io_out_kv(local_pes_16_7_io_out_kv),
    .io_out_stage(local_pes_16_7_io_out_stage)
  );
  PE_1 local_pes_16_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_8_clock),
    .reset(local_pes_16_8_reset),
    .io_in_q(local_pes_16_8_io_in_q),
    .io_in_sum(local_pes_16_8_io_in_sum),
    .io_in_sum_exp(local_pes_16_8_io_in_sum_exp),
    .io_in_kv(local_pes_16_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_8_io_in_inv_sum),
    .io_in_stage(local_pes_16_8_io_in_stage),
    .io_out_q(local_pes_16_8_io_out_q),
    .io_out_sum(local_pes_16_8_io_out_sum),
    .io_out_sum_exp(local_pes_16_8_io_out_sum_exp),
    .io_out_kv(local_pes_16_8_io_out_kv),
    .io_out_stage(local_pes_16_8_io_out_stage)
  );
  PE_1 local_pes_16_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_9_clock),
    .reset(local_pes_16_9_reset),
    .io_in_q(local_pes_16_9_io_in_q),
    .io_in_sum(local_pes_16_9_io_in_sum),
    .io_in_sum_exp(local_pes_16_9_io_in_sum_exp),
    .io_in_kv(local_pes_16_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_9_io_in_inv_sum),
    .io_in_stage(local_pes_16_9_io_in_stage),
    .io_out_q(local_pes_16_9_io_out_q),
    .io_out_sum(local_pes_16_9_io_out_sum),
    .io_out_sum_exp(local_pes_16_9_io_out_sum_exp),
    .io_out_kv(local_pes_16_9_io_out_kv),
    .io_out_stage(local_pes_16_9_io_out_stage)
  );
  PE_1 local_pes_16_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_10_clock),
    .reset(local_pes_16_10_reset),
    .io_in_q(local_pes_16_10_io_in_q),
    .io_in_sum(local_pes_16_10_io_in_sum),
    .io_in_sum_exp(local_pes_16_10_io_in_sum_exp),
    .io_in_kv(local_pes_16_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_10_io_in_inv_sum),
    .io_in_stage(local_pes_16_10_io_in_stage),
    .io_out_q(local_pes_16_10_io_out_q),
    .io_out_sum(local_pes_16_10_io_out_sum),
    .io_out_sum_exp(local_pes_16_10_io_out_sum_exp),
    .io_out_kv(local_pes_16_10_io_out_kv),
    .io_out_stage(local_pes_16_10_io_out_stage)
  );
  PE_1 local_pes_16_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_11_clock),
    .reset(local_pes_16_11_reset),
    .io_in_q(local_pes_16_11_io_in_q),
    .io_in_sum(local_pes_16_11_io_in_sum),
    .io_in_sum_exp(local_pes_16_11_io_in_sum_exp),
    .io_in_kv(local_pes_16_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_11_io_in_inv_sum),
    .io_in_stage(local_pes_16_11_io_in_stage),
    .io_out_q(local_pes_16_11_io_out_q),
    .io_out_sum(local_pes_16_11_io_out_sum),
    .io_out_sum_exp(local_pes_16_11_io_out_sum_exp),
    .io_out_kv(local_pes_16_11_io_out_kv),
    .io_out_stage(local_pes_16_11_io_out_stage)
  );
  PE_1 local_pes_16_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_12_clock),
    .reset(local_pes_16_12_reset),
    .io_in_q(local_pes_16_12_io_in_q),
    .io_in_sum(local_pes_16_12_io_in_sum),
    .io_in_sum_exp(local_pes_16_12_io_in_sum_exp),
    .io_in_kv(local_pes_16_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_12_io_in_inv_sum),
    .io_in_stage(local_pes_16_12_io_in_stage),
    .io_out_q(local_pes_16_12_io_out_q),
    .io_out_sum(local_pes_16_12_io_out_sum),
    .io_out_sum_exp(local_pes_16_12_io_out_sum_exp),
    .io_out_kv(local_pes_16_12_io_out_kv),
    .io_out_stage(local_pes_16_12_io_out_stage)
  );
  PE_1 local_pes_16_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_13_clock),
    .reset(local_pes_16_13_reset),
    .io_in_q(local_pes_16_13_io_in_q),
    .io_in_sum(local_pes_16_13_io_in_sum),
    .io_in_sum_exp(local_pes_16_13_io_in_sum_exp),
    .io_in_kv(local_pes_16_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_13_io_in_inv_sum),
    .io_in_stage(local_pes_16_13_io_in_stage),
    .io_out_q(local_pes_16_13_io_out_q),
    .io_out_sum(local_pes_16_13_io_out_sum),
    .io_out_sum_exp(local_pes_16_13_io_out_sum_exp),
    .io_out_kv(local_pes_16_13_io_out_kv),
    .io_out_stage(local_pes_16_13_io_out_stage)
  );
  PE_1 local_pes_16_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_14_clock),
    .reset(local_pes_16_14_reset),
    .io_in_q(local_pes_16_14_io_in_q),
    .io_in_sum(local_pes_16_14_io_in_sum),
    .io_in_sum_exp(local_pes_16_14_io_in_sum_exp),
    .io_in_kv(local_pes_16_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_14_io_in_inv_sum),
    .io_in_stage(local_pes_16_14_io_in_stage),
    .io_out_q(local_pes_16_14_io_out_q),
    .io_out_sum(local_pes_16_14_io_out_sum),
    .io_out_sum_exp(local_pes_16_14_io_out_sum_exp),
    .io_out_kv(local_pes_16_14_io_out_kv),
    .io_out_stage(local_pes_16_14_io_out_stage)
  );
  PE_1 local_pes_16_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_15_clock),
    .reset(local_pes_16_15_reset),
    .io_in_q(local_pes_16_15_io_in_q),
    .io_in_sum(local_pes_16_15_io_in_sum),
    .io_in_sum_exp(local_pes_16_15_io_in_sum_exp),
    .io_in_kv(local_pes_16_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_15_io_in_inv_sum),
    .io_in_stage(local_pes_16_15_io_in_stage),
    .io_out_q(local_pes_16_15_io_out_q),
    .io_out_sum(local_pes_16_15_io_out_sum),
    .io_out_sum_exp(local_pes_16_15_io_out_sum_exp),
    .io_out_kv(local_pes_16_15_io_out_kv),
    .io_out_stage(local_pes_16_15_io_out_stage)
  );
  PE_1 local_pes_16_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_16_clock),
    .reset(local_pes_16_16_reset),
    .io_in_q(local_pes_16_16_io_in_q),
    .io_in_sum(local_pes_16_16_io_in_sum),
    .io_in_sum_exp(local_pes_16_16_io_in_sum_exp),
    .io_in_kv(local_pes_16_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_16_io_in_inv_sum),
    .io_in_stage(local_pes_16_16_io_in_stage),
    .io_out_q(local_pes_16_16_io_out_q),
    .io_out_sum(local_pes_16_16_io_out_sum),
    .io_out_sum_exp(local_pes_16_16_io_out_sum_exp),
    .io_out_kv(local_pes_16_16_io_out_kv),
    .io_out_stage(local_pes_16_16_io_out_stage)
  );
  PE_1 local_pes_16_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_17_clock),
    .reset(local_pes_16_17_reset),
    .io_in_q(local_pes_16_17_io_in_q),
    .io_in_sum(local_pes_16_17_io_in_sum),
    .io_in_sum_exp(local_pes_16_17_io_in_sum_exp),
    .io_in_kv(local_pes_16_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_17_io_in_inv_sum),
    .io_in_stage(local_pes_16_17_io_in_stage),
    .io_out_q(local_pes_16_17_io_out_q),
    .io_out_sum(local_pes_16_17_io_out_sum),
    .io_out_sum_exp(local_pes_16_17_io_out_sum_exp),
    .io_out_kv(local_pes_16_17_io_out_kv),
    .io_out_stage(local_pes_16_17_io_out_stage)
  );
  PE_1 local_pes_16_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_18_clock),
    .reset(local_pes_16_18_reset),
    .io_in_q(local_pes_16_18_io_in_q),
    .io_in_sum(local_pes_16_18_io_in_sum),
    .io_in_sum_exp(local_pes_16_18_io_in_sum_exp),
    .io_in_kv(local_pes_16_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_18_io_in_inv_sum),
    .io_in_stage(local_pes_16_18_io_in_stage),
    .io_out_q(local_pes_16_18_io_out_q),
    .io_out_sum(local_pes_16_18_io_out_sum),
    .io_out_sum_exp(local_pes_16_18_io_out_sum_exp),
    .io_out_kv(local_pes_16_18_io_out_kv),
    .io_out_stage(local_pes_16_18_io_out_stage)
  );
  PE_1 local_pes_16_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_19_clock),
    .reset(local_pes_16_19_reset),
    .io_in_q(local_pes_16_19_io_in_q),
    .io_in_sum(local_pes_16_19_io_in_sum),
    .io_in_sum_exp(local_pes_16_19_io_in_sum_exp),
    .io_in_kv(local_pes_16_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_19_io_in_inv_sum),
    .io_in_stage(local_pes_16_19_io_in_stage),
    .io_out_q(local_pes_16_19_io_out_q),
    .io_out_sum(local_pes_16_19_io_out_sum),
    .io_out_sum_exp(local_pes_16_19_io_out_sum_exp),
    .io_out_kv(local_pes_16_19_io_out_kv),
    .io_out_stage(local_pes_16_19_io_out_stage)
  );
  PE_1 local_pes_16_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_20_clock),
    .reset(local_pes_16_20_reset),
    .io_in_q(local_pes_16_20_io_in_q),
    .io_in_sum(local_pes_16_20_io_in_sum),
    .io_in_sum_exp(local_pes_16_20_io_in_sum_exp),
    .io_in_kv(local_pes_16_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_20_io_in_inv_sum),
    .io_in_stage(local_pes_16_20_io_in_stage),
    .io_out_q(local_pes_16_20_io_out_q),
    .io_out_sum(local_pes_16_20_io_out_sum),
    .io_out_sum_exp(local_pes_16_20_io_out_sum_exp),
    .io_out_kv(local_pes_16_20_io_out_kv),
    .io_out_stage(local_pes_16_20_io_out_stage)
  );
  PE_1 local_pes_16_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_21_clock),
    .reset(local_pes_16_21_reset),
    .io_in_q(local_pes_16_21_io_in_q),
    .io_in_sum(local_pes_16_21_io_in_sum),
    .io_in_sum_exp(local_pes_16_21_io_in_sum_exp),
    .io_in_kv(local_pes_16_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_21_io_in_inv_sum),
    .io_in_stage(local_pes_16_21_io_in_stage),
    .io_out_q(local_pes_16_21_io_out_q),
    .io_out_sum(local_pes_16_21_io_out_sum),
    .io_out_sum_exp(local_pes_16_21_io_out_sum_exp),
    .io_out_kv(local_pes_16_21_io_out_kv),
    .io_out_stage(local_pes_16_21_io_out_stage)
  );
  PE_1 local_pes_16_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_22_clock),
    .reset(local_pes_16_22_reset),
    .io_in_q(local_pes_16_22_io_in_q),
    .io_in_sum(local_pes_16_22_io_in_sum),
    .io_in_sum_exp(local_pes_16_22_io_in_sum_exp),
    .io_in_kv(local_pes_16_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_22_io_in_inv_sum),
    .io_in_stage(local_pes_16_22_io_in_stage),
    .io_out_q(local_pes_16_22_io_out_q),
    .io_out_sum(local_pes_16_22_io_out_sum),
    .io_out_sum_exp(local_pes_16_22_io_out_sum_exp),
    .io_out_kv(local_pes_16_22_io_out_kv),
    .io_out_stage(local_pes_16_22_io_out_stage)
  );
  PE_1 local_pes_16_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_23_clock),
    .reset(local_pes_16_23_reset),
    .io_in_q(local_pes_16_23_io_in_q),
    .io_in_sum(local_pes_16_23_io_in_sum),
    .io_in_sum_exp(local_pes_16_23_io_in_sum_exp),
    .io_in_kv(local_pes_16_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_23_io_in_inv_sum),
    .io_in_stage(local_pes_16_23_io_in_stage),
    .io_out_q(local_pes_16_23_io_out_q),
    .io_out_sum(local_pes_16_23_io_out_sum),
    .io_out_sum_exp(local_pes_16_23_io_out_sum_exp),
    .io_out_kv(local_pes_16_23_io_out_kv),
    .io_out_stage(local_pes_16_23_io_out_stage)
  );
  PE_1 local_pes_16_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_24_clock),
    .reset(local_pes_16_24_reset),
    .io_in_q(local_pes_16_24_io_in_q),
    .io_in_sum(local_pes_16_24_io_in_sum),
    .io_in_sum_exp(local_pes_16_24_io_in_sum_exp),
    .io_in_kv(local_pes_16_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_24_io_in_inv_sum),
    .io_in_stage(local_pes_16_24_io_in_stage),
    .io_out_q(local_pes_16_24_io_out_q),
    .io_out_sum(local_pes_16_24_io_out_sum),
    .io_out_sum_exp(local_pes_16_24_io_out_sum_exp),
    .io_out_kv(local_pes_16_24_io_out_kv),
    .io_out_stage(local_pes_16_24_io_out_stage)
  );
  PE_1 local_pes_16_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_25_clock),
    .reset(local_pes_16_25_reset),
    .io_in_q(local_pes_16_25_io_in_q),
    .io_in_sum(local_pes_16_25_io_in_sum),
    .io_in_sum_exp(local_pes_16_25_io_in_sum_exp),
    .io_in_kv(local_pes_16_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_25_io_in_inv_sum),
    .io_in_stage(local_pes_16_25_io_in_stage),
    .io_out_q(local_pes_16_25_io_out_q),
    .io_out_sum(local_pes_16_25_io_out_sum),
    .io_out_sum_exp(local_pes_16_25_io_out_sum_exp),
    .io_out_kv(local_pes_16_25_io_out_kv),
    .io_out_stage(local_pes_16_25_io_out_stage)
  );
  PE_1 local_pes_16_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_26_clock),
    .reset(local_pes_16_26_reset),
    .io_in_q(local_pes_16_26_io_in_q),
    .io_in_sum(local_pes_16_26_io_in_sum),
    .io_in_sum_exp(local_pes_16_26_io_in_sum_exp),
    .io_in_kv(local_pes_16_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_26_io_in_inv_sum),
    .io_in_stage(local_pes_16_26_io_in_stage),
    .io_out_q(local_pes_16_26_io_out_q),
    .io_out_sum(local_pes_16_26_io_out_sum),
    .io_out_sum_exp(local_pes_16_26_io_out_sum_exp),
    .io_out_kv(local_pes_16_26_io_out_kv),
    .io_out_stage(local_pes_16_26_io_out_stage)
  );
  PE_1 local_pes_16_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_27_clock),
    .reset(local_pes_16_27_reset),
    .io_in_q(local_pes_16_27_io_in_q),
    .io_in_sum(local_pes_16_27_io_in_sum),
    .io_in_sum_exp(local_pes_16_27_io_in_sum_exp),
    .io_in_kv(local_pes_16_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_27_io_in_inv_sum),
    .io_in_stage(local_pes_16_27_io_in_stage),
    .io_out_q(local_pes_16_27_io_out_q),
    .io_out_sum(local_pes_16_27_io_out_sum),
    .io_out_sum_exp(local_pes_16_27_io_out_sum_exp),
    .io_out_kv(local_pes_16_27_io_out_kv),
    .io_out_stage(local_pes_16_27_io_out_stage)
  );
  PE_1 local_pes_16_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_28_clock),
    .reset(local_pes_16_28_reset),
    .io_in_q(local_pes_16_28_io_in_q),
    .io_in_sum(local_pes_16_28_io_in_sum),
    .io_in_sum_exp(local_pes_16_28_io_in_sum_exp),
    .io_in_kv(local_pes_16_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_28_io_in_inv_sum),
    .io_in_stage(local_pes_16_28_io_in_stage),
    .io_out_q(local_pes_16_28_io_out_q),
    .io_out_sum(local_pes_16_28_io_out_sum),
    .io_out_sum_exp(local_pes_16_28_io_out_sum_exp),
    .io_out_kv(local_pes_16_28_io_out_kv),
    .io_out_stage(local_pes_16_28_io_out_stage)
  );
  PE_1 local_pes_16_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_29_clock),
    .reset(local_pes_16_29_reset),
    .io_in_q(local_pes_16_29_io_in_q),
    .io_in_sum(local_pes_16_29_io_in_sum),
    .io_in_sum_exp(local_pes_16_29_io_in_sum_exp),
    .io_in_kv(local_pes_16_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_29_io_in_inv_sum),
    .io_in_stage(local_pes_16_29_io_in_stage),
    .io_out_q(local_pes_16_29_io_out_q),
    .io_out_sum(local_pes_16_29_io_out_sum),
    .io_out_sum_exp(local_pes_16_29_io_out_sum_exp),
    .io_out_kv(local_pes_16_29_io_out_kv),
    .io_out_stage(local_pes_16_29_io_out_stage)
  );
  PE_1 local_pes_16_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_30_clock),
    .reset(local_pes_16_30_reset),
    .io_in_q(local_pes_16_30_io_in_q),
    .io_in_sum(local_pes_16_30_io_in_sum),
    .io_in_sum_exp(local_pes_16_30_io_in_sum_exp),
    .io_in_kv(local_pes_16_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_30_io_in_inv_sum),
    .io_in_stage(local_pes_16_30_io_in_stage),
    .io_out_q(local_pes_16_30_io_out_q),
    .io_out_sum(local_pes_16_30_io_out_sum),
    .io_out_sum_exp(local_pes_16_30_io_out_sum_exp),
    .io_out_kv(local_pes_16_30_io_out_kv),
    .io_out_stage(local_pes_16_30_io_out_stage)
  );
  PE_1 local_pes_16_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_16_31_clock),
    .reset(local_pes_16_31_reset),
    .io_in_q(local_pes_16_31_io_in_q),
    .io_in_sum(local_pes_16_31_io_in_sum),
    .io_in_sum_exp(local_pes_16_31_io_in_sum_exp),
    .io_in_kv(local_pes_16_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_16_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_16_31_io_in_inv_sum),
    .io_in_stage(local_pes_16_31_io_in_stage),
    .io_out_q(local_pes_16_31_io_out_q),
    .io_out_sum(local_pes_16_31_io_out_sum),
    .io_out_sum_exp(local_pes_16_31_io_out_sum_exp),
    .io_out_kv(local_pes_16_31_io_out_kv),
    .io_out_stage(local_pes_16_31_io_out_stage)
  );
  PE local_pes_17_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_0_clock),
    .reset(local_pes_17_0_reset),
    .io_in_q(local_pes_17_0_io_in_q),
    .io_in_kv(local_pes_17_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_0_io_in_inv_sum),
    .io_in_stage(local_pes_17_0_io_in_stage),
    .io_out_q(local_pes_17_0_io_out_q),
    .io_out_sum(local_pes_17_0_io_out_sum),
    .io_out_kv(local_pes_17_0_io_out_kv),
    .io_out_stage(local_pes_17_0_io_out_stage)
  );
  PE_1 local_pes_17_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_1_clock),
    .reset(local_pes_17_1_reset),
    .io_in_q(local_pes_17_1_io_in_q),
    .io_in_sum(local_pes_17_1_io_in_sum),
    .io_in_sum_exp(local_pes_17_1_io_in_sum_exp),
    .io_in_kv(local_pes_17_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_1_io_in_inv_sum),
    .io_in_stage(local_pes_17_1_io_in_stage),
    .io_out_q(local_pes_17_1_io_out_q),
    .io_out_sum(local_pes_17_1_io_out_sum),
    .io_out_sum_exp(local_pes_17_1_io_out_sum_exp),
    .io_out_kv(local_pes_17_1_io_out_kv),
    .io_out_stage(local_pes_17_1_io_out_stage)
  );
  PE_1 local_pes_17_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_2_clock),
    .reset(local_pes_17_2_reset),
    .io_in_q(local_pes_17_2_io_in_q),
    .io_in_sum(local_pes_17_2_io_in_sum),
    .io_in_sum_exp(local_pes_17_2_io_in_sum_exp),
    .io_in_kv(local_pes_17_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_2_io_in_inv_sum),
    .io_in_stage(local_pes_17_2_io_in_stage),
    .io_out_q(local_pes_17_2_io_out_q),
    .io_out_sum(local_pes_17_2_io_out_sum),
    .io_out_sum_exp(local_pes_17_2_io_out_sum_exp),
    .io_out_kv(local_pes_17_2_io_out_kv),
    .io_out_stage(local_pes_17_2_io_out_stage)
  );
  PE_1 local_pes_17_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_3_clock),
    .reset(local_pes_17_3_reset),
    .io_in_q(local_pes_17_3_io_in_q),
    .io_in_sum(local_pes_17_3_io_in_sum),
    .io_in_sum_exp(local_pes_17_3_io_in_sum_exp),
    .io_in_kv(local_pes_17_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_3_io_in_inv_sum),
    .io_in_stage(local_pes_17_3_io_in_stage),
    .io_out_q(local_pes_17_3_io_out_q),
    .io_out_sum(local_pes_17_3_io_out_sum),
    .io_out_sum_exp(local_pes_17_3_io_out_sum_exp),
    .io_out_kv(local_pes_17_3_io_out_kv),
    .io_out_stage(local_pes_17_3_io_out_stage)
  );
  PE_1 local_pes_17_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_4_clock),
    .reset(local_pes_17_4_reset),
    .io_in_q(local_pes_17_4_io_in_q),
    .io_in_sum(local_pes_17_4_io_in_sum),
    .io_in_sum_exp(local_pes_17_4_io_in_sum_exp),
    .io_in_kv(local_pes_17_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_4_io_in_inv_sum),
    .io_in_stage(local_pes_17_4_io_in_stage),
    .io_out_q(local_pes_17_4_io_out_q),
    .io_out_sum(local_pes_17_4_io_out_sum),
    .io_out_sum_exp(local_pes_17_4_io_out_sum_exp),
    .io_out_kv(local_pes_17_4_io_out_kv),
    .io_out_stage(local_pes_17_4_io_out_stage)
  );
  PE_1 local_pes_17_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_5_clock),
    .reset(local_pes_17_5_reset),
    .io_in_q(local_pes_17_5_io_in_q),
    .io_in_sum(local_pes_17_5_io_in_sum),
    .io_in_sum_exp(local_pes_17_5_io_in_sum_exp),
    .io_in_kv(local_pes_17_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_5_io_in_inv_sum),
    .io_in_stage(local_pes_17_5_io_in_stage),
    .io_out_q(local_pes_17_5_io_out_q),
    .io_out_sum(local_pes_17_5_io_out_sum),
    .io_out_sum_exp(local_pes_17_5_io_out_sum_exp),
    .io_out_kv(local_pes_17_5_io_out_kv),
    .io_out_stage(local_pes_17_5_io_out_stage)
  );
  PE_1 local_pes_17_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_6_clock),
    .reset(local_pes_17_6_reset),
    .io_in_q(local_pes_17_6_io_in_q),
    .io_in_sum(local_pes_17_6_io_in_sum),
    .io_in_sum_exp(local_pes_17_6_io_in_sum_exp),
    .io_in_kv(local_pes_17_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_6_io_in_inv_sum),
    .io_in_stage(local_pes_17_6_io_in_stage),
    .io_out_q(local_pes_17_6_io_out_q),
    .io_out_sum(local_pes_17_6_io_out_sum),
    .io_out_sum_exp(local_pes_17_6_io_out_sum_exp),
    .io_out_kv(local_pes_17_6_io_out_kv),
    .io_out_stage(local_pes_17_6_io_out_stage)
  );
  PE_1 local_pes_17_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_7_clock),
    .reset(local_pes_17_7_reset),
    .io_in_q(local_pes_17_7_io_in_q),
    .io_in_sum(local_pes_17_7_io_in_sum),
    .io_in_sum_exp(local_pes_17_7_io_in_sum_exp),
    .io_in_kv(local_pes_17_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_7_io_in_inv_sum),
    .io_in_stage(local_pes_17_7_io_in_stage),
    .io_out_q(local_pes_17_7_io_out_q),
    .io_out_sum(local_pes_17_7_io_out_sum),
    .io_out_sum_exp(local_pes_17_7_io_out_sum_exp),
    .io_out_kv(local_pes_17_7_io_out_kv),
    .io_out_stage(local_pes_17_7_io_out_stage)
  );
  PE_1 local_pes_17_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_8_clock),
    .reset(local_pes_17_8_reset),
    .io_in_q(local_pes_17_8_io_in_q),
    .io_in_sum(local_pes_17_8_io_in_sum),
    .io_in_sum_exp(local_pes_17_8_io_in_sum_exp),
    .io_in_kv(local_pes_17_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_8_io_in_inv_sum),
    .io_in_stage(local_pes_17_8_io_in_stage),
    .io_out_q(local_pes_17_8_io_out_q),
    .io_out_sum(local_pes_17_8_io_out_sum),
    .io_out_sum_exp(local_pes_17_8_io_out_sum_exp),
    .io_out_kv(local_pes_17_8_io_out_kv),
    .io_out_stage(local_pes_17_8_io_out_stage)
  );
  PE_1 local_pes_17_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_9_clock),
    .reset(local_pes_17_9_reset),
    .io_in_q(local_pes_17_9_io_in_q),
    .io_in_sum(local_pes_17_9_io_in_sum),
    .io_in_sum_exp(local_pes_17_9_io_in_sum_exp),
    .io_in_kv(local_pes_17_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_9_io_in_inv_sum),
    .io_in_stage(local_pes_17_9_io_in_stage),
    .io_out_q(local_pes_17_9_io_out_q),
    .io_out_sum(local_pes_17_9_io_out_sum),
    .io_out_sum_exp(local_pes_17_9_io_out_sum_exp),
    .io_out_kv(local_pes_17_9_io_out_kv),
    .io_out_stage(local_pes_17_9_io_out_stage)
  );
  PE_1 local_pes_17_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_10_clock),
    .reset(local_pes_17_10_reset),
    .io_in_q(local_pes_17_10_io_in_q),
    .io_in_sum(local_pes_17_10_io_in_sum),
    .io_in_sum_exp(local_pes_17_10_io_in_sum_exp),
    .io_in_kv(local_pes_17_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_10_io_in_inv_sum),
    .io_in_stage(local_pes_17_10_io_in_stage),
    .io_out_q(local_pes_17_10_io_out_q),
    .io_out_sum(local_pes_17_10_io_out_sum),
    .io_out_sum_exp(local_pes_17_10_io_out_sum_exp),
    .io_out_kv(local_pes_17_10_io_out_kv),
    .io_out_stage(local_pes_17_10_io_out_stage)
  );
  PE_1 local_pes_17_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_11_clock),
    .reset(local_pes_17_11_reset),
    .io_in_q(local_pes_17_11_io_in_q),
    .io_in_sum(local_pes_17_11_io_in_sum),
    .io_in_sum_exp(local_pes_17_11_io_in_sum_exp),
    .io_in_kv(local_pes_17_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_11_io_in_inv_sum),
    .io_in_stage(local_pes_17_11_io_in_stage),
    .io_out_q(local_pes_17_11_io_out_q),
    .io_out_sum(local_pes_17_11_io_out_sum),
    .io_out_sum_exp(local_pes_17_11_io_out_sum_exp),
    .io_out_kv(local_pes_17_11_io_out_kv),
    .io_out_stage(local_pes_17_11_io_out_stage)
  );
  PE_1 local_pes_17_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_12_clock),
    .reset(local_pes_17_12_reset),
    .io_in_q(local_pes_17_12_io_in_q),
    .io_in_sum(local_pes_17_12_io_in_sum),
    .io_in_sum_exp(local_pes_17_12_io_in_sum_exp),
    .io_in_kv(local_pes_17_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_12_io_in_inv_sum),
    .io_in_stage(local_pes_17_12_io_in_stage),
    .io_out_q(local_pes_17_12_io_out_q),
    .io_out_sum(local_pes_17_12_io_out_sum),
    .io_out_sum_exp(local_pes_17_12_io_out_sum_exp),
    .io_out_kv(local_pes_17_12_io_out_kv),
    .io_out_stage(local_pes_17_12_io_out_stage)
  );
  PE_1 local_pes_17_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_13_clock),
    .reset(local_pes_17_13_reset),
    .io_in_q(local_pes_17_13_io_in_q),
    .io_in_sum(local_pes_17_13_io_in_sum),
    .io_in_sum_exp(local_pes_17_13_io_in_sum_exp),
    .io_in_kv(local_pes_17_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_13_io_in_inv_sum),
    .io_in_stage(local_pes_17_13_io_in_stage),
    .io_out_q(local_pes_17_13_io_out_q),
    .io_out_sum(local_pes_17_13_io_out_sum),
    .io_out_sum_exp(local_pes_17_13_io_out_sum_exp),
    .io_out_kv(local_pes_17_13_io_out_kv),
    .io_out_stage(local_pes_17_13_io_out_stage)
  );
  PE_1 local_pes_17_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_14_clock),
    .reset(local_pes_17_14_reset),
    .io_in_q(local_pes_17_14_io_in_q),
    .io_in_sum(local_pes_17_14_io_in_sum),
    .io_in_sum_exp(local_pes_17_14_io_in_sum_exp),
    .io_in_kv(local_pes_17_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_14_io_in_inv_sum),
    .io_in_stage(local_pes_17_14_io_in_stage),
    .io_out_q(local_pes_17_14_io_out_q),
    .io_out_sum(local_pes_17_14_io_out_sum),
    .io_out_sum_exp(local_pes_17_14_io_out_sum_exp),
    .io_out_kv(local_pes_17_14_io_out_kv),
    .io_out_stage(local_pes_17_14_io_out_stage)
  );
  PE_1 local_pes_17_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_15_clock),
    .reset(local_pes_17_15_reset),
    .io_in_q(local_pes_17_15_io_in_q),
    .io_in_sum(local_pes_17_15_io_in_sum),
    .io_in_sum_exp(local_pes_17_15_io_in_sum_exp),
    .io_in_kv(local_pes_17_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_15_io_in_inv_sum),
    .io_in_stage(local_pes_17_15_io_in_stage),
    .io_out_q(local_pes_17_15_io_out_q),
    .io_out_sum(local_pes_17_15_io_out_sum),
    .io_out_sum_exp(local_pes_17_15_io_out_sum_exp),
    .io_out_kv(local_pes_17_15_io_out_kv),
    .io_out_stage(local_pes_17_15_io_out_stage)
  );
  PE_1 local_pes_17_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_16_clock),
    .reset(local_pes_17_16_reset),
    .io_in_q(local_pes_17_16_io_in_q),
    .io_in_sum(local_pes_17_16_io_in_sum),
    .io_in_sum_exp(local_pes_17_16_io_in_sum_exp),
    .io_in_kv(local_pes_17_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_16_io_in_inv_sum),
    .io_in_stage(local_pes_17_16_io_in_stage),
    .io_out_q(local_pes_17_16_io_out_q),
    .io_out_sum(local_pes_17_16_io_out_sum),
    .io_out_sum_exp(local_pes_17_16_io_out_sum_exp),
    .io_out_kv(local_pes_17_16_io_out_kv),
    .io_out_stage(local_pes_17_16_io_out_stage)
  );
  PE_1 local_pes_17_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_17_clock),
    .reset(local_pes_17_17_reset),
    .io_in_q(local_pes_17_17_io_in_q),
    .io_in_sum(local_pes_17_17_io_in_sum),
    .io_in_sum_exp(local_pes_17_17_io_in_sum_exp),
    .io_in_kv(local_pes_17_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_17_io_in_inv_sum),
    .io_in_stage(local_pes_17_17_io_in_stage),
    .io_out_q(local_pes_17_17_io_out_q),
    .io_out_sum(local_pes_17_17_io_out_sum),
    .io_out_sum_exp(local_pes_17_17_io_out_sum_exp),
    .io_out_kv(local_pes_17_17_io_out_kv),
    .io_out_stage(local_pes_17_17_io_out_stage)
  );
  PE_1 local_pes_17_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_18_clock),
    .reset(local_pes_17_18_reset),
    .io_in_q(local_pes_17_18_io_in_q),
    .io_in_sum(local_pes_17_18_io_in_sum),
    .io_in_sum_exp(local_pes_17_18_io_in_sum_exp),
    .io_in_kv(local_pes_17_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_18_io_in_inv_sum),
    .io_in_stage(local_pes_17_18_io_in_stage),
    .io_out_q(local_pes_17_18_io_out_q),
    .io_out_sum(local_pes_17_18_io_out_sum),
    .io_out_sum_exp(local_pes_17_18_io_out_sum_exp),
    .io_out_kv(local_pes_17_18_io_out_kv),
    .io_out_stage(local_pes_17_18_io_out_stage)
  );
  PE_1 local_pes_17_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_19_clock),
    .reset(local_pes_17_19_reset),
    .io_in_q(local_pes_17_19_io_in_q),
    .io_in_sum(local_pes_17_19_io_in_sum),
    .io_in_sum_exp(local_pes_17_19_io_in_sum_exp),
    .io_in_kv(local_pes_17_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_19_io_in_inv_sum),
    .io_in_stage(local_pes_17_19_io_in_stage),
    .io_out_q(local_pes_17_19_io_out_q),
    .io_out_sum(local_pes_17_19_io_out_sum),
    .io_out_sum_exp(local_pes_17_19_io_out_sum_exp),
    .io_out_kv(local_pes_17_19_io_out_kv),
    .io_out_stage(local_pes_17_19_io_out_stage)
  );
  PE_1 local_pes_17_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_20_clock),
    .reset(local_pes_17_20_reset),
    .io_in_q(local_pes_17_20_io_in_q),
    .io_in_sum(local_pes_17_20_io_in_sum),
    .io_in_sum_exp(local_pes_17_20_io_in_sum_exp),
    .io_in_kv(local_pes_17_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_20_io_in_inv_sum),
    .io_in_stage(local_pes_17_20_io_in_stage),
    .io_out_q(local_pes_17_20_io_out_q),
    .io_out_sum(local_pes_17_20_io_out_sum),
    .io_out_sum_exp(local_pes_17_20_io_out_sum_exp),
    .io_out_kv(local_pes_17_20_io_out_kv),
    .io_out_stage(local_pes_17_20_io_out_stage)
  );
  PE_1 local_pes_17_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_21_clock),
    .reset(local_pes_17_21_reset),
    .io_in_q(local_pes_17_21_io_in_q),
    .io_in_sum(local_pes_17_21_io_in_sum),
    .io_in_sum_exp(local_pes_17_21_io_in_sum_exp),
    .io_in_kv(local_pes_17_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_21_io_in_inv_sum),
    .io_in_stage(local_pes_17_21_io_in_stage),
    .io_out_q(local_pes_17_21_io_out_q),
    .io_out_sum(local_pes_17_21_io_out_sum),
    .io_out_sum_exp(local_pes_17_21_io_out_sum_exp),
    .io_out_kv(local_pes_17_21_io_out_kv),
    .io_out_stage(local_pes_17_21_io_out_stage)
  );
  PE_1 local_pes_17_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_22_clock),
    .reset(local_pes_17_22_reset),
    .io_in_q(local_pes_17_22_io_in_q),
    .io_in_sum(local_pes_17_22_io_in_sum),
    .io_in_sum_exp(local_pes_17_22_io_in_sum_exp),
    .io_in_kv(local_pes_17_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_22_io_in_inv_sum),
    .io_in_stage(local_pes_17_22_io_in_stage),
    .io_out_q(local_pes_17_22_io_out_q),
    .io_out_sum(local_pes_17_22_io_out_sum),
    .io_out_sum_exp(local_pes_17_22_io_out_sum_exp),
    .io_out_kv(local_pes_17_22_io_out_kv),
    .io_out_stage(local_pes_17_22_io_out_stage)
  );
  PE_1 local_pes_17_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_23_clock),
    .reset(local_pes_17_23_reset),
    .io_in_q(local_pes_17_23_io_in_q),
    .io_in_sum(local_pes_17_23_io_in_sum),
    .io_in_sum_exp(local_pes_17_23_io_in_sum_exp),
    .io_in_kv(local_pes_17_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_23_io_in_inv_sum),
    .io_in_stage(local_pes_17_23_io_in_stage),
    .io_out_q(local_pes_17_23_io_out_q),
    .io_out_sum(local_pes_17_23_io_out_sum),
    .io_out_sum_exp(local_pes_17_23_io_out_sum_exp),
    .io_out_kv(local_pes_17_23_io_out_kv),
    .io_out_stage(local_pes_17_23_io_out_stage)
  );
  PE_1 local_pes_17_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_24_clock),
    .reset(local_pes_17_24_reset),
    .io_in_q(local_pes_17_24_io_in_q),
    .io_in_sum(local_pes_17_24_io_in_sum),
    .io_in_sum_exp(local_pes_17_24_io_in_sum_exp),
    .io_in_kv(local_pes_17_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_24_io_in_inv_sum),
    .io_in_stage(local_pes_17_24_io_in_stage),
    .io_out_q(local_pes_17_24_io_out_q),
    .io_out_sum(local_pes_17_24_io_out_sum),
    .io_out_sum_exp(local_pes_17_24_io_out_sum_exp),
    .io_out_kv(local_pes_17_24_io_out_kv),
    .io_out_stage(local_pes_17_24_io_out_stage)
  );
  PE_1 local_pes_17_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_25_clock),
    .reset(local_pes_17_25_reset),
    .io_in_q(local_pes_17_25_io_in_q),
    .io_in_sum(local_pes_17_25_io_in_sum),
    .io_in_sum_exp(local_pes_17_25_io_in_sum_exp),
    .io_in_kv(local_pes_17_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_25_io_in_inv_sum),
    .io_in_stage(local_pes_17_25_io_in_stage),
    .io_out_q(local_pes_17_25_io_out_q),
    .io_out_sum(local_pes_17_25_io_out_sum),
    .io_out_sum_exp(local_pes_17_25_io_out_sum_exp),
    .io_out_kv(local_pes_17_25_io_out_kv),
    .io_out_stage(local_pes_17_25_io_out_stage)
  );
  PE_1 local_pes_17_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_26_clock),
    .reset(local_pes_17_26_reset),
    .io_in_q(local_pes_17_26_io_in_q),
    .io_in_sum(local_pes_17_26_io_in_sum),
    .io_in_sum_exp(local_pes_17_26_io_in_sum_exp),
    .io_in_kv(local_pes_17_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_26_io_in_inv_sum),
    .io_in_stage(local_pes_17_26_io_in_stage),
    .io_out_q(local_pes_17_26_io_out_q),
    .io_out_sum(local_pes_17_26_io_out_sum),
    .io_out_sum_exp(local_pes_17_26_io_out_sum_exp),
    .io_out_kv(local_pes_17_26_io_out_kv),
    .io_out_stage(local_pes_17_26_io_out_stage)
  );
  PE_1 local_pes_17_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_27_clock),
    .reset(local_pes_17_27_reset),
    .io_in_q(local_pes_17_27_io_in_q),
    .io_in_sum(local_pes_17_27_io_in_sum),
    .io_in_sum_exp(local_pes_17_27_io_in_sum_exp),
    .io_in_kv(local_pes_17_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_27_io_in_inv_sum),
    .io_in_stage(local_pes_17_27_io_in_stage),
    .io_out_q(local_pes_17_27_io_out_q),
    .io_out_sum(local_pes_17_27_io_out_sum),
    .io_out_sum_exp(local_pes_17_27_io_out_sum_exp),
    .io_out_kv(local_pes_17_27_io_out_kv),
    .io_out_stage(local_pes_17_27_io_out_stage)
  );
  PE_1 local_pes_17_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_28_clock),
    .reset(local_pes_17_28_reset),
    .io_in_q(local_pes_17_28_io_in_q),
    .io_in_sum(local_pes_17_28_io_in_sum),
    .io_in_sum_exp(local_pes_17_28_io_in_sum_exp),
    .io_in_kv(local_pes_17_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_28_io_in_inv_sum),
    .io_in_stage(local_pes_17_28_io_in_stage),
    .io_out_q(local_pes_17_28_io_out_q),
    .io_out_sum(local_pes_17_28_io_out_sum),
    .io_out_sum_exp(local_pes_17_28_io_out_sum_exp),
    .io_out_kv(local_pes_17_28_io_out_kv),
    .io_out_stage(local_pes_17_28_io_out_stage)
  );
  PE_1 local_pes_17_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_29_clock),
    .reset(local_pes_17_29_reset),
    .io_in_q(local_pes_17_29_io_in_q),
    .io_in_sum(local_pes_17_29_io_in_sum),
    .io_in_sum_exp(local_pes_17_29_io_in_sum_exp),
    .io_in_kv(local_pes_17_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_29_io_in_inv_sum),
    .io_in_stage(local_pes_17_29_io_in_stage),
    .io_out_q(local_pes_17_29_io_out_q),
    .io_out_sum(local_pes_17_29_io_out_sum),
    .io_out_sum_exp(local_pes_17_29_io_out_sum_exp),
    .io_out_kv(local_pes_17_29_io_out_kv),
    .io_out_stage(local_pes_17_29_io_out_stage)
  );
  PE_1 local_pes_17_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_30_clock),
    .reset(local_pes_17_30_reset),
    .io_in_q(local_pes_17_30_io_in_q),
    .io_in_sum(local_pes_17_30_io_in_sum),
    .io_in_sum_exp(local_pes_17_30_io_in_sum_exp),
    .io_in_kv(local_pes_17_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_30_io_in_inv_sum),
    .io_in_stage(local_pes_17_30_io_in_stage),
    .io_out_q(local_pes_17_30_io_out_q),
    .io_out_sum(local_pes_17_30_io_out_sum),
    .io_out_sum_exp(local_pes_17_30_io_out_sum_exp),
    .io_out_kv(local_pes_17_30_io_out_kv),
    .io_out_stage(local_pes_17_30_io_out_stage)
  );
  PE_1 local_pes_17_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_17_31_clock),
    .reset(local_pes_17_31_reset),
    .io_in_q(local_pes_17_31_io_in_q),
    .io_in_sum(local_pes_17_31_io_in_sum),
    .io_in_sum_exp(local_pes_17_31_io_in_sum_exp),
    .io_in_kv(local_pes_17_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_17_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_17_31_io_in_inv_sum),
    .io_in_stage(local_pes_17_31_io_in_stage),
    .io_out_q(local_pes_17_31_io_out_q),
    .io_out_sum(local_pes_17_31_io_out_sum),
    .io_out_sum_exp(local_pes_17_31_io_out_sum_exp),
    .io_out_kv(local_pes_17_31_io_out_kv),
    .io_out_stage(local_pes_17_31_io_out_stage)
  );
  PE local_pes_18_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_0_clock),
    .reset(local_pes_18_0_reset),
    .io_in_q(local_pes_18_0_io_in_q),
    .io_in_kv(local_pes_18_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_0_io_in_inv_sum),
    .io_in_stage(local_pes_18_0_io_in_stage),
    .io_out_q(local_pes_18_0_io_out_q),
    .io_out_sum(local_pes_18_0_io_out_sum),
    .io_out_kv(local_pes_18_0_io_out_kv),
    .io_out_stage(local_pes_18_0_io_out_stage)
  );
  PE_1 local_pes_18_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_1_clock),
    .reset(local_pes_18_1_reset),
    .io_in_q(local_pes_18_1_io_in_q),
    .io_in_sum(local_pes_18_1_io_in_sum),
    .io_in_sum_exp(local_pes_18_1_io_in_sum_exp),
    .io_in_kv(local_pes_18_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_1_io_in_inv_sum),
    .io_in_stage(local_pes_18_1_io_in_stage),
    .io_out_q(local_pes_18_1_io_out_q),
    .io_out_sum(local_pes_18_1_io_out_sum),
    .io_out_sum_exp(local_pes_18_1_io_out_sum_exp),
    .io_out_kv(local_pes_18_1_io_out_kv),
    .io_out_stage(local_pes_18_1_io_out_stage)
  );
  PE_1 local_pes_18_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_2_clock),
    .reset(local_pes_18_2_reset),
    .io_in_q(local_pes_18_2_io_in_q),
    .io_in_sum(local_pes_18_2_io_in_sum),
    .io_in_sum_exp(local_pes_18_2_io_in_sum_exp),
    .io_in_kv(local_pes_18_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_2_io_in_inv_sum),
    .io_in_stage(local_pes_18_2_io_in_stage),
    .io_out_q(local_pes_18_2_io_out_q),
    .io_out_sum(local_pes_18_2_io_out_sum),
    .io_out_sum_exp(local_pes_18_2_io_out_sum_exp),
    .io_out_kv(local_pes_18_2_io_out_kv),
    .io_out_stage(local_pes_18_2_io_out_stage)
  );
  PE_1 local_pes_18_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_3_clock),
    .reset(local_pes_18_3_reset),
    .io_in_q(local_pes_18_3_io_in_q),
    .io_in_sum(local_pes_18_3_io_in_sum),
    .io_in_sum_exp(local_pes_18_3_io_in_sum_exp),
    .io_in_kv(local_pes_18_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_3_io_in_inv_sum),
    .io_in_stage(local_pes_18_3_io_in_stage),
    .io_out_q(local_pes_18_3_io_out_q),
    .io_out_sum(local_pes_18_3_io_out_sum),
    .io_out_sum_exp(local_pes_18_3_io_out_sum_exp),
    .io_out_kv(local_pes_18_3_io_out_kv),
    .io_out_stage(local_pes_18_3_io_out_stage)
  );
  PE_1 local_pes_18_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_4_clock),
    .reset(local_pes_18_4_reset),
    .io_in_q(local_pes_18_4_io_in_q),
    .io_in_sum(local_pes_18_4_io_in_sum),
    .io_in_sum_exp(local_pes_18_4_io_in_sum_exp),
    .io_in_kv(local_pes_18_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_4_io_in_inv_sum),
    .io_in_stage(local_pes_18_4_io_in_stage),
    .io_out_q(local_pes_18_4_io_out_q),
    .io_out_sum(local_pes_18_4_io_out_sum),
    .io_out_sum_exp(local_pes_18_4_io_out_sum_exp),
    .io_out_kv(local_pes_18_4_io_out_kv),
    .io_out_stage(local_pes_18_4_io_out_stage)
  );
  PE_1 local_pes_18_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_5_clock),
    .reset(local_pes_18_5_reset),
    .io_in_q(local_pes_18_5_io_in_q),
    .io_in_sum(local_pes_18_5_io_in_sum),
    .io_in_sum_exp(local_pes_18_5_io_in_sum_exp),
    .io_in_kv(local_pes_18_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_5_io_in_inv_sum),
    .io_in_stage(local_pes_18_5_io_in_stage),
    .io_out_q(local_pes_18_5_io_out_q),
    .io_out_sum(local_pes_18_5_io_out_sum),
    .io_out_sum_exp(local_pes_18_5_io_out_sum_exp),
    .io_out_kv(local_pes_18_5_io_out_kv),
    .io_out_stage(local_pes_18_5_io_out_stage)
  );
  PE_1 local_pes_18_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_6_clock),
    .reset(local_pes_18_6_reset),
    .io_in_q(local_pes_18_6_io_in_q),
    .io_in_sum(local_pes_18_6_io_in_sum),
    .io_in_sum_exp(local_pes_18_6_io_in_sum_exp),
    .io_in_kv(local_pes_18_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_6_io_in_inv_sum),
    .io_in_stage(local_pes_18_6_io_in_stage),
    .io_out_q(local_pes_18_6_io_out_q),
    .io_out_sum(local_pes_18_6_io_out_sum),
    .io_out_sum_exp(local_pes_18_6_io_out_sum_exp),
    .io_out_kv(local_pes_18_6_io_out_kv),
    .io_out_stage(local_pes_18_6_io_out_stage)
  );
  PE_1 local_pes_18_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_7_clock),
    .reset(local_pes_18_7_reset),
    .io_in_q(local_pes_18_7_io_in_q),
    .io_in_sum(local_pes_18_7_io_in_sum),
    .io_in_sum_exp(local_pes_18_7_io_in_sum_exp),
    .io_in_kv(local_pes_18_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_7_io_in_inv_sum),
    .io_in_stage(local_pes_18_7_io_in_stage),
    .io_out_q(local_pes_18_7_io_out_q),
    .io_out_sum(local_pes_18_7_io_out_sum),
    .io_out_sum_exp(local_pes_18_7_io_out_sum_exp),
    .io_out_kv(local_pes_18_7_io_out_kv),
    .io_out_stage(local_pes_18_7_io_out_stage)
  );
  PE_1 local_pes_18_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_8_clock),
    .reset(local_pes_18_8_reset),
    .io_in_q(local_pes_18_8_io_in_q),
    .io_in_sum(local_pes_18_8_io_in_sum),
    .io_in_sum_exp(local_pes_18_8_io_in_sum_exp),
    .io_in_kv(local_pes_18_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_8_io_in_inv_sum),
    .io_in_stage(local_pes_18_8_io_in_stage),
    .io_out_q(local_pes_18_8_io_out_q),
    .io_out_sum(local_pes_18_8_io_out_sum),
    .io_out_sum_exp(local_pes_18_8_io_out_sum_exp),
    .io_out_kv(local_pes_18_8_io_out_kv),
    .io_out_stage(local_pes_18_8_io_out_stage)
  );
  PE_1 local_pes_18_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_9_clock),
    .reset(local_pes_18_9_reset),
    .io_in_q(local_pes_18_9_io_in_q),
    .io_in_sum(local_pes_18_9_io_in_sum),
    .io_in_sum_exp(local_pes_18_9_io_in_sum_exp),
    .io_in_kv(local_pes_18_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_9_io_in_inv_sum),
    .io_in_stage(local_pes_18_9_io_in_stage),
    .io_out_q(local_pes_18_9_io_out_q),
    .io_out_sum(local_pes_18_9_io_out_sum),
    .io_out_sum_exp(local_pes_18_9_io_out_sum_exp),
    .io_out_kv(local_pes_18_9_io_out_kv),
    .io_out_stage(local_pes_18_9_io_out_stage)
  );
  PE_1 local_pes_18_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_10_clock),
    .reset(local_pes_18_10_reset),
    .io_in_q(local_pes_18_10_io_in_q),
    .io_in_sum(local_pes_18_10_io_in_sum),
    .io_in_sum_exp(local_pes_18_10_io_in_sum_exp),
    .io_in_kv(local_pes_18_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_10_io_in_inv_sum),
    .io_in_stage(local_pes_18_10_io_in_stage),
    .io_out_q(local_pes_18_10_io_out_q),
    .io_out_sum(local_pes_18_10_io_out_sum),
    .io_out_sum_exp(local_pes_18_10_io_out_sum_exp),
    .io_out_kv(local_pes_18_10_io_out_kv),
    .io_out_stage(local_pes_18_10_io_out_stage)
  );
  PE_1 local_pes_18_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_11_clock),
    .reset(local_pes_18_11_reset),
    .io_in_q(local_pes_18_11_io_in_q),
    .io_in_sum(local_pes_18_11_io_in_sum),
    .io_in_sum_exp(local_pes_18_11_io_in_sum_exp),
    .io_in_kv(local_pes_18_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_11_io_in_inv_sum),
    .io_in_stage(local_pes_18_11_io_in_stage),
    .io_out_q(local_pes_18_11_io_out_q),
    .io_out_sum(local_pes_18_11_io_out_sum),
    .io_out_sum_exp(local_pes_18_11_io_out_sum_exp),
    .io_out_kv(local_pes_18_11_io_out_kv),
    .io_out_stage(local_pes_18_11_io_out_stage)
  );
  PE_1 local_pes_18_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_12_clock),
    .reset(local_pes_18_12_reset),
    .io_in_q(local_pes_18_12_io_in_q),
    .io_in_sum(local_pes_18_12_io_in_sum),
    .io_in_sum_exp(local_pes_18_12_io_in_sum_exp),
    .io_in_kv(local_pes_18_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_12_io_in_inv_sum),
    .io_in_stage(local_pes_18_12_io_in_stage),
    .io_out_q(local_pes_18_12_io_out_q),
    .io_out_sum(local_pes_18_12_io_out_sum),
    .io_out_sum_exp(local_pes_18_12_io_out_sum_exp),
    .io_out_kv(local_pes_18_12_io_out_kv),
    .io_out_stage(local_pes_18_12_io_out_stage)
  );
  PE_1 local_pes_18_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_13_clock),
    .reset(local_pes_18_13_reset),
    .io_in_q(local_pes_18_13_io_in_q),
    .io_in_sum(local_pes_18_13_io_in_sum),
    .io_in_sum_exp(local_pes_18_13_io_in_sum_exp),
    .io_in_kv(local_pes_18_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_13_io_in_inv_sum),
    .io_in_stage(local_pes_18_13_io_in_stage),
    .io_out_q(local_pes_18_13_io_out_q),
    .io_out_sum(local_pes_18_13_io_out_sum),
    .io_out_sum_exp(local_pes_18_13_io_out_sum_exp),
    .io_out_kv(local_pes_18_13_io_out_kv),
    .io_out_stage(local_pes_18_13_io_out_stage)
  );
  PE_1 local_pes_18_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_14_clock),
    .reset(local_pes_18_14_reset),
    .io_in_q(local_pes_18_14_io_in_q),
    .io_in_sum(local_pes_18_14_io_in_sum),
    .io_in_sum_exp(local_pes_18_14_io_in_sum_exp),
    .io_in_kv(local_pes_18_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_14_io_in_inv_sum),
    .io_in_stage(local_pes_18_14_io_in_stage),
    .io_out_q(local_pes_18_14_io_out_q),
    .io_out_sum(local_pes_18_14_io_out_sum),
    .io_out_sum_exp(local_pes_18_14_io_out_sum_exp),
    .io_out_kv(local_pes_18_14_io_out_kv),
    .io_out_stage(local_pes_18_14_io_out_stage)
  );
  PE_1 local_pes_18_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_15_clock),
    .reset(local_pes_18_15_reset),
    .io_in_q(local_pes_18_15_io_in_q),
    .io_in_sum(local_pes_18_15_io_in_sum),
    .io_in_sum_exp(local_pes_18_15_io_in_sum_exp),
    .io_in_kv(local_pes_18_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_15_io_in_inv_sum),
    .io_in_stage(local_pes_18_15_io_in_stage),
    .io_out_q(local_pes_18_15_io_out_q),
    .io_out_sum(local_pes_18_15_io_out_sum),
    .io_out_sum_exp(local_pes_18_15_io_out_sum_exp),
    .io_out_kv(local_pes_18_15_io_out_kv),
    .io_out_stage(local_pes_18_15_io_out_stage)
  );
  PE_1 local_pes_18_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_16_clock),
    .reset(local_pes_18_16_reset),
    .io_in_q(local_pes_18_16_io_in_q),
    .io_in_sum(local_pes_18_16_io_in_sum),
    .io_in_sum_exp(local_pes_18_16_io_in_sum_exp),
    .io_in_kv(local_pes_18_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_16_io_in_inv_sum),
    .io_in_stage(local_pes_18_16_io_in_stage),
    .io_out_q(local_pes_18_16_io_out_q),
    .io_out_sum(local_pes_18_16_io_out_sum),
    .io_out_sum_exp(local_pes_18_16_io_out_sum_exp),
    .io_out_kv(local_pes_18_16_io_out_kv),
    .io_out_stage(local_pes_18_16_io_out_stage)
  );
  PE_1 local_pes_18_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_17_clock),
    .reset(local_pes_18_17_reset),
    .io_in_q(local_pes_18_17_io_in_q),
    .io_in_sum(local_pes_18_17_io_in_sum),
    .io_in_sum_exp(local_pes_18_17_io_in_sum_exp),
    .io_in_kv(local_pes_18_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_17_io_in_inv_sum),
    .io_in_stage(local_pes_18_17_io_in_stage),
    .io_out_q(local_pes_18_17_io_out_q),
    .io_out_sum(local_pes_18_17_io_out_sum),
    .io_out_sum_exp(local_pes_18_17_io_out_sum_exp),
    .io_out_kv(local_pes_18_17_io_out_kv),
    .io_out_stage(local_pes_18_17_io_out_stage)
  );
  PE_1 local_pes_18_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_18_clock),
    .reset(local_pes_18_18_reset),
    .io_in_q(local_pes_18_18_io_in_q),
    .io_in_sum(local_pes_18_18_io_in_sum),
    .io_in_sum_exp(local_pes_18_18_io_in_sum_exp),
    .io_in_kv(local_pes_18_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_18_io_in_inv_sum),
    .io_in_stage(local_pes_18_18_io_in_stage),
    .io_out_q(local_pes_18_18_io_out_q),
    .io_out_sum(local_pes_18_18_io_out_sum),
    .io_out_sum_exp(local_pes_18_18_io_out_sum_exp),
    .io_out_kv(local_pes_18_18_io_out_kv),
    .io_out_stage(local_pes_18_18_io_out_stage)
  );
  PE_1 local_pes_18_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_19_clock),
    .reset(local_pes_18_19_reset),
    .io_in_q(local_pes_18_19_io_in_q),
    .io_in_sum(local_pes_18_19_io_in_sum),
    .io_in_sum_exp(local_pes_18_19_io_in_sum_exp),
    .io_in_kv(local_pes_18_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_19_io_in_inv_sum),
    .io_in_stage(local_pes_18_19_io_in_stage),
    .io_out_q(local_pes_18_19_io_out_q),
    .io_out_sum(local_pes_18_19_io_out_sum),
    .io_out_sum_exp(local_pes_18_19_io_out_sum_exp),
    .io_out_kv(local_pes_18_19_io_out_kv),
    .io_out_stage(local_pes_18_19_io_out_stage)
  );
  PE_1 local_pes_18_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_20_clock),
    .reset(local_pes_18_20_reset),
    .io_in_q(local_pes_18_20_io_in_q),
    .io_in_sum(local_pes_18_20_io_in_sum),
    .io_in_sum_exp(local_pes_18_20_io_in_sum_exp),
    .io_in_kv(local_pes_18_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_20_io_in_inv_sum),
    .io_in_stage(local_pes_18_20_io_in_stage),
    .io_out_q(local_pes_18_20_io_out_q),
    .io_out_sum(local_pes_18_20_io_out_sum),
    .io_out_sum_exp(local_pes_18_20_io_out_sum_exp),
    .io_out_kv(local_pes_18_20_io_out_kv),
    .io_out_stage(local_pes_18_20_io_out_stage)
  );
  PE_1 local_pes_18_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_21_clock),
    .reset(local_pes_18_21_reset),
    .io_in_q(local_pes_18_21_io_in_q),
    .io_in_sum(local_pes_18_21_io_in_sum),
    .io_in_sum_exp(local_pes_18_21_io_in_sum_exp),
    .io_in_kv(local_pes_18_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_21_io_in_inv_sum),
    .io_in_stage(local_pes_18_21_io_in_stage),
    .io_out_q(local_pes_18_21_io_out_q),
    .io_out_sum(local_pes_18_21_io_out_sum),
    .io_out_sum_exp(local_pes_18_21_io_out_sum_exp),
    .io_out_kv(local_pes_18_21_io_out_kv),
    .io_out_stage(local_pes_18_21_io_out_stage)
  );
  PE_1 local_pes_18_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_22_clock),
    .reset(local_pes_18_22_reset),
    .io_in_q(local_pes_18_22_io_in_q),
    .io_in_sum(local_pes_18_22_io_in_sum),
    .io_in_sum_exp(local_pes_18_22_io_in_sum_exp),
    .io_in_kv(local_pes_18_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_22_io_in_inv_sum),
    .io_in_stage(local_pes_18_22_io_in_stage),
    .io_out_q(local_pes_18_22_io_out_q),
    .io_out_sum(local_pes_18_22_io_out_sum),
    .io_out_sum_exp(local_pes_18_22_io_out_sum_exp),
    .io_out_kv(local_pes_18_22_io_out_kv),
    .io_out_stage(local_pes_18_22_io_out_stage)
  );
  PE_1 local_pes_18_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_23_clock),
    .reset(local_pes_18_23_reset),
    .io_in_q(local_pes_18_23_io_in_q),
    .io_in_sum(local_pes_18_23_io_in_sum),
    .io_in_sum_exp(local_pes_18_23_io_in_sum_exp),
    .io_in_kv(local_pes_18_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_23_io_in_inv_sum),
    .io_in_stage(local_pes_18_23_io_in_stage),
    .io_out_q(local_pes_18_23_io_out_q),
    .io_out_sum(local_pes_18_23_io_out_sum),
    .io_out_sum_exp(local_pes_18_23_io_out_sum_exp),
    .io_out_kv(local_pes_18_23_io_out_kv),
    .io_out_stage(local_pes_18_23_io_out_stage)
  );
  PE_1 local_pes_18_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_24_clock),
    .reset(local_pes_18_24_reset),
    .io_in_q(local_pes_18_24_io_in_q),
    .io_in_sum(local_pes_18_24_io_in_sum),
    .io_in_sum_exp(local_pes_18_24_io_in_sum_exp),
    .io_in_kv(local_pes_18_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_24_io_in_inv_sum),
    .io_in_stage(local_pes_18_24_io_in_stage),
    .io_out_q(local_pes_18_24_io_out_q),
    .io_out_sum(local_pes_18_24_io_out_sum),
    .io_out_sum_exp(local_pes_18_24_io_out_sum_exp),
    .io_out_kv(local_pes_18_24_io_out_kv),
    .io_out_stage(local_pes_18_24_io_out_stage)
  );
  PE_1 local_pes_18_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_25_clock),
    .reset(local_pes_18_25_reset),
    .io_in_q(local_pes_18_25_io_in_q),
    .io_in_sum(local_pes_18_25_io_in_sum),
    .io_in_sum_exp(local_pes_18_25_io_in_sum_exp),
    .io_in_kv(local_pes_18_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_25_io_in_inv_sum),
    .io_in_stage(local_pes_18_25_io_in_stage),
    .io_out_q(local_pes_18_25_io_out_q),
    .io_out_sum(local_pes_18_25_io_out_sum),
    .io_out_sum_exp(local_pes_18_25_io_out_sum_exp),
    .io_out_kv(local_pes_18_25_io_out_kv),
    .io_out_stage(local_pes_18_25_io_out_stage)
  );
  PE_1 local_pes_18_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_26_clock),
    .reset(local_pes_18_26_reset),
    .io_in_q(local_pes_18_26_io_in_q),
    .io_in_sum(local_pes_18_26_io_in_sum),
    .io_in_sum_exp(local_pes_18_26_io_in_sum_exp),
    .io_in_kv(local_pes_18_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_26_io_in_inv_sum),
    .io_in_stage(local_pes_18_26_io_in_stage),
    .io_out_q(local_pes_18_26_io_out_q),
    .io_out_sum(local_pes_18_26_io_out_sum),
    .io_out_sum_exp(local_pes_18_26_io_out_sum_exp),
    .io_out_kv(local_pes_18_26_io_out_kv),
    .io_out_stage(local_pes_18_26_io_out_stage)
  );
  PE_1 local_pes_18_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_27_clock),
    .reset(local_pes_18_27_reset),
    .io_in_q(local_pes_18_27_io_in_q),
    .io_in_sum(local_pes_18_27_io_in_sum),
    .io_in_sum_exp(local_pes_18_27_io_in_sum_exp),
    .io_in_kv(local_pes_18_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_27_io_in_inv_sum),
    .io_in_stage(local_pes_18_27_io_in_stage),
    .io_out_q(local_pes_18_27_io_out_q),
    .io_out_sum(local_pes_18_27_io_out_sum),
    .io_out_sum_exp(local_pes_18_27_io_out_sum_exp),
    .io_out_kv(local_pes_18_27_io_out_kv),
    .io_out_stage(local_pes_18_27_io_out_stage)
  );
  PE_1 local_pes_18_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_28_clock),
    .reset(local_pes_18_28_reset),
    .io_in_q(local_pes_18_28_io_in_q),
    .io_in_sum(local_pes_18_28_io_in_sum),
    .io_in_sum_exp(local_pes_18_28_io_in_sum_exp),
    .io_in_kv(local_pes_18_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_28_io_in_inv_sum),
    .io_in_stage(local_pes_18_28_io_in_stage),
    .io_out_q(local_pes_18_28_io_out_q),
    .io_out_sum(local_pes_18_28_io_out_sum),
    .io_out_sum_exp(local_pes_18_28_io_out_sum_exp),
    .io_out_kv(local_pes_18_28_io_out_kv),
    .io_out_stage(local_pes_18_28_io_out_stage)
  );
  PE_1 local_pes_18_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_29_clock),
    .reset(local_pes_18_29_reset),
    .io_in_q(local_pes_18_29_io_in_q),
    .io_in_sum(local_pes_18_29_io_in_sum),
    .io_in_sum_exp(local_pes_18_29_io_in_sum_exp),
    .io_in_kv(local_pes_18_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_29_io_in_inv_sum),
    .io_in_stage(local_pes_18_29_io_in_stage),
    .io_out_q(local_pes_18_29_io_out_q),
    .io_out_sum(local_pes_18_29_io_out_sum),
    .io_out_sum_exp(local_pes_18_29_io_out_sum_exp),
    .io_out_kv(local_pes_18_29_io_out_kv),
    .io_out_stage(local_pes_18_29_io_out_stage)
  );
  PE_1 local_pes_18_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_30_clock),
    .reset(local_pes_18_30_reset),
    .io_in_q(local_pes_18_30_io_in_q),
    .io_in_sum(local_pes_18_30_io_in_sum),
    .io_in_sum_exp(local_pes_18_30_io_in_sum_exp),
    .io_in_kv(local_pes_18_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_30_io_in_inv_sum),
    .io_in_stage(local_pes_18_30_io_in_stage),
    .io_out_q(local_pes_18_30_io_out_q),
    .io_out_sum(local_pes_18_30_io_out_sum),
    .io_out_sum_exp(local_pes_18_30_io_out_sum_exp),
    .io_out_kv(local_pes_18_30_io_out_kv),
    .io_out_stage(local_pes_18_30_io_out_stage)
  );
  PE_1 local_pes_18_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_18_31_clock),
    .reset(local_pes_18_31_reset),
    .io_in_q(local_pes_18_31_io_in_q),
    .io_in_sum(local_pes_18_31_io_in_sum),
    .io_in_sum_exp(local_pes_18_31_io_in_sum_exp),
    .io_in_kv(local_pes_18_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_18_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_18_31_io_in_inv_sum),
    .io_in_stage(local_pes_18_31_io_in_stage),
    .io_out_q(local_pes_18_31_io_out_q),
    .io_out_sum(local_pes_18_31_io_out_sum),
    .io_out_sum_exp(local_pes_18_31_io_out_sum_exp),
    .io_out_kv(local_pes_18_31_io_out_kv),
    .io_out_stage(local_pes_18_31_io_out_stage)
  );
  PE local_pes_19_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_0_clock),
    .reset(local_pes_19_0_reset),
    .io_in_q(local_pes_19_0_io_in_q),
    .io_in_kv(local_pes_19_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_0_io_in_inv_sum),
    .io_in_stage(local_pes_19_0_io_in_stage),
    .io_out_q(local_pes_19_0_io_out_q),
    .io_out_sum(local_pes_19_0_io_out_sum),
    .io_out_kv(local_pes_19_0_io_out_kv),
    .io_out_stage(local_pes_19_0_io_out_stage)
  );
  PE_1 local_pes_19_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_1_clock),
    .reset(local_pes_19_1_reset),
    .io_in_q(local_pes_19_1_io_in_q),
    .io_in_sum(local_pes_19_1_io_in_sum),
    .io_in_sum_exp(local_pes_19_1_io_in_sum_exp),
    .io_in_kv(local_pes_19_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_1_io_in_inv_sum),
    .io_in_stage(local_pes_19_1_io_in_stage),
    .io_out_q(local_pes_19_1_io_out_q),
    .io_out_sum(local_pes_19_1_io_out_sum),
    .io_out_sum_exp(local_pes_19_1_io_out_sum_exp),
    .io_out_kv(local_pes_19_1_io_out_kv),
    .io_out_stage(local_pes_19_1_io_out_stage)
  );
  PE_1 local_pes_19_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_2_clock),
    .reset(local_pes_19_2_reset),
    .io_in_q(local_pes_19_2_io_in_q),
    .io_in_sum(local_pes_19_2_io_in_sum),
    .io_in_sum_exp(local_pes_19_2_io_in_sum_exp),
    .io_in_kv(local_pes_19_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_2_io_in_inv_sum),
    .io_in_stage(local_pes_19_2_io_in_stage),
    .io_out_q(local_pes_19_2_io_out_q),
    .io_out_sum(local_pes_19_2_io_out_sum),
    .io_out_sum_exp(local_pes_19_2_io_out_sum_exp),
    .io_out_kv(local_pes_19_2_io_out_kv),
    .io_out_stage(local_pes_19_2_io_out_stage)
  );
  PE_1 local_pes_19_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_3_clock),
    .reset(local_pes_19_3_reset),
    .io_in_q(local_pes_19_3_io_in_q),
    .io_in_sum(local_pes_19_3_io_in_sum),
    .io_in_sum_exp(local_pes_19_3_io_in_sum_exp),
    .io_in_kv(local_pes_19_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_3_io_in_inv_sum),
    .io_in_stage(local_pes_19_3_io_in_stage),
    .io_out_q(local_pes_19_3_io_out_q),
    .io_out_sum(local_pes_19_3_io_out_sum),
    .io_out_sum_exp(local_pes_19_3_io_out_sum_exp),
    .io_out_kv(local_pes_19_3_io_out_kv),
    .io_out_stage(local_pes_19_3_io_out_stage)
  );
  PE_1 local_pes_19_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_4_clock),
    .reset(local_pes_19_4_reset),
    .io_in_q(local_pes_19_4_io_in_q),
    .io_in_sum(local_pes_19_4_io_in_sum),
    .io_in_sum_exp(local_pes_19_4_io_in_sum_exp),
    .io_in_kv(local_pes_19_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_4_io_in_inv_sum),
    .io_in_stage(local_pes_19_4_io_in_stage),
    .io_out_q(local_pes_19_4_io_out_q),
    .io_out_sum(local_pes_19_4_io_out_sum),
    .io_out_sum_exp(local_pes_19_4_io_out_sum_exp),
    .io_out_kv(local_pes_19_4_io_out_kv),
    .io_out_stage(local_pes_19_4_io_out_stage)
  );
  PE_1 local_pes_19_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_5_clock),
    .reset(local_pes_19_5_reset),
    .io_in_q(local_pes_19_5_io_in_q),
    .io_in_sum(local_pes_19_5_io_in_sum),
    .io_in_sum_exp(local_pes_19_5_io_in_sum_exp),
    .io_in_kv(local_pes_19_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_5_io_in_inv_sum),
    .io_in_stage(local_pes_19_5_io_in_stage),
    .io_out_q(local_pes_19_5_io_out_q),
    .io_out_sum(local_pes_19_5_io_out_sum),
    .io_out_sum_exp(local_pes_19_5_io_out_sum_exp),
    .io_out_kv(local_pes_19_5_io_out_kv),
    .io_out_stage(local_pes_19_5_io_out_stage)
  );
  PE_1 local_pes_19_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_6_clock),
    .reset(local_pes_19_6_reset),
    .io_in_q(local_pes_19_6_io_in_q),
    .io_in_sum(local_pes_19_6_io_in_sum),
    .io_in_sum_exp(local_pes_19_6_io_in_sum_exp),
    .io_in_kv(local_pes_19_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_6_io_in_inv_sum),
    .io_in_stage(local_pes_19_6_io_in_stage),
    .io_out_q(local_pes_19_6_io_out_q),
    .io_out_sum(local_pes_19_6_io_out_sum),
    .io_out_sum_exp(local_pes_19_6_io_out_sum_exp),
    .io_out_kv(local_pes_19_6_io_out_kv),
    .io_out_stage(local_pes_19_6_io_out_stage)
  );
  PE_1 local_pes_19_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_7_clock),
    .reset(local_pes_19_7_reset),
    .io_in_q(local_pes_19_7_io_in_q),
    .io_in_sum(local_pes_19_7_io_in_sum),
    .io_in_sum_exp(local_pes_19_7_io_in_sum_exp),
    .io_in_kv(local_pes_19_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_7_io_in_inv_sum),
    .io_in_stage(local_pes_19_7_io_in_stage),
    .io_out_q(local_pes_19_7_io_out_q),
    .io_out_sum(local_pes_19_7_io_out_sum),
    .io_out_sum_exp(local_pes_19_7_io_out_sum_exp),
    .io_out_kv(local_pes_19_7_io_out_kv),
    .io_out_stage(local_pes_19_7_io_out_stage)
  );
  PE_1 local_pes_19_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_8_clock),
    .reset(local_pes_19_8_reset),
    .io_in_q(local_pes_19_8_io_in_q),
    .io_in_sum(local_pes_19_8_io_in_sum),
    .io_in_sum_exp(local_pes_19_8_io_in_sum_exp),
    .io_in_kv(local_pes_19_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_8_io_in_inv_sum),
    .io_in_stage(local_pes_19_8_io_in_stage),
    .io_out_q(local_pes_19_8_io_out_q),
    .io_out_sum(local_pes_19_8_io_out_sum),
    .io_out_sum_exp(local_pes_19_8_io_out_sum_exp),
    .io_out_kv(local_pes_19_8_io_out_kv),
    .io_out_stage(local_pes_19_8_io_out_stage)
  );
  PE_1 local_pes_19_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_9_clock),
    .reset(local_pes_19_9_reset),
    .io_in_q(local_pes_19_9_io_in_q),
    .io_in_sum(local_pes_19_9_io_in_sum),
    .io_in_sum_exp(local_pes_19_9_io_in_sum_exp),
    .io_in_kv(local_pes_19_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_9_io_in_inv_sum),
    .io_in_stage(local_pes_19_9_io_in_stage),
    .io_out_q(local_pes_19_9_io_out_q),
    .io_out_sum(local_pes_19_9_io_out_sum),
    .io_out_sum_exp(local_pes_19_9_io_out_sum_exp),
    .io_out_kv(local_pes_19_9_io_out_kv),
    .io_out_stage(local_pes_19_9_io_out_stage)
  );
  PE_1 local_pes_19_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_10_clock),
    .reset(local_pes_19_10_reset),
    .io_in_q(local_pes_19_10_io_in_q),
    .io_in_sum(local_pes_19_10_io_in_sum),
    .io_in_sum_exp(local_pes_19_10_io_in_sum_exp),
    .io_in_kv(local_pes_19_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_10_io_in_inv_sum),
    .io_in_stage(local_pes_19_10_io_in_stage),
    .io_out_q(local_pes_19_10_io_out_q),
    .io_out_sum(local_pes_19_10_io_out_sum),
    .io_out_sum_exp(local_pes_19_10_io_out_sum_exp),
    .io_out_kv(local_pes_19_10_io_out_kv),
    .io_out_stage(local_pes_19_10_io_out_stage)
  );
  PE_1 local_pes_19_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_11_clock),
    .reset(local_pes_19_11_reset),
    .io_in_q(local_pes_19_11_io_in_q),
    .io_in_sum(local_pes_19_11_io_in_sum),
    .io_in_sum_exp(local_pes_19_11_io_in_sum_exp),
    .io_in_kv(local_pes_19_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_11_io_in_inv_sum),
    .io_in_stage(local_pes_19_11_io_in_stage),
    .io_out_q(local_pes_19_11_io_out_q),
    .io_out_sum(local_pes_19_11_io_out_sum),
    .io_out_sum_exp(local_pes_19_11_io_out_sum_exp),
    .io_out_kv(local_pes_19_11_io_out_kv),
    .io_out_stage(local_pes_19_11_io_out_stage)
  );
  PE_1 local_pes_19_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_12_clock),
    .reset(local_pes_19_12_reset),
    .io_in_q(local_pes_19_12_io_in_q),
    .io_in_sum(local_pes_19_12_io_in_sum),
    .io_in_sum_exp(local_pes_19_12_io_in_sum_exp),
    .io_in_kv(local_pes_19_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_12_io_in_inv_sum),
    .io_in_stage(local_pes_19_12_io_in_stage),
    .io_out_q(local_pes_19_12_io_out_q),
    .io_out_sum(local_pes_19_12_io_out_sum),
    .io_out_sum_exp(local_pes_19_12_io_out_sum_exp),
    .io_out_kv(local_pes_19_12_io_out_kv),
    .io_out_stage(local_pes_19_12_io_out_stage)
  );
  PE_1 local_pes_19_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_13_clock),
    .reset(local_pes_19_13_reset),
    .io_in_q(local_pes_19_13_io_in_q),
    .io_in_sum(local_pes_19_13_io_in_sum),
    .io_in_sum_exp(local_pes_19_13_io_in_sum_exp),
    .io_in_kv(local_pes_19_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_13_io_in_inv_sum),
    .io_in_stage(local_pes_19_13_io_in_stage),
    .io_out_q(local_pes_19_13_io_out_q),
    .io_out_sum(local_pes_19_13_io_out_sum),
    .io_out_sum_exp(local_pes_19_13_io_out_sum_exp),
    .io_out_kv(local_pes_19_13_io_out_kv),
    .io_out_stage(local_pes_19_13_io_out_stage)
  );
  PE_1 local_pes_19_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_14_clock),
    .reset(local_pes_19_14_reset),
    .io_in_q(local_pes_19_14_io_in_q),
    .io_in_sum(local_pes_19_14_io_in_sum),
    .io_in_sum_exp(local_pes_19_14_io_in_sum_exp),
    .io_in_kv(local_pes_19_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_14_io_in_inv_sum),
    .io_in_stage(local_pes_19_14_io_in_stage),
    .io_out_q(local_pes_19_14_io_out_q),
    .io_out_sum(local_pes_19_14_io_out_sum),
    .io_out_sum_exp(local_pes_19_14_io_out_sum_exp),
    .io_out_kv(local_pes_19_14_io_out_kv),
    .io_out_stage(local_pes_19_14_io_out_stage)
  );
  PE_1 local_pes_19_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_15_clock),
    .reset(local_pes_19_15_reset),
    .io_in_q(local_pes_19_15_io_in_q),
    .io_in_sum(local_pes_19_15_io_in_sum),
    .io_in_sum_exp(local_pes_19_15_io_in_sum_exp),
    .io_in_kv(local_pes_19_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_15_io_in_inv_sum),
    .io_in_stage(local_pes_19_15_io_in_stage),
    .io_out_q(local_pes_19_15_io_out_q),
    .io_out_sum(local_pes_19_15_io_out_sum),
    .io_out_sum_exp(local_pes_19_15_io_out_sum_exp),
    .io_out_kv(local_pes_19_15_io_out_kv),
    .io_out_stage(local_pes_19_15_io_out_stage)
  );
  PE_1 local_pes_19_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_16_clock),
    .reset(local_pes_19_16_reset),
    .io_in_q(local_pes_19_16_io_in_q),
    .io_in_sum(local_pes_19_16_io_in_sum),
    .io_in_sum_exp(local_pes_19_16_io_in_sum_exp),
    .io_in_kv(local_pes_19_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_16_io_in_inv_sum),
    .io_in_stage(local_pes_19_16_io_in_stage),
    .io_out_q(local_pes_19_16_io_out_q),
    .io_out_sum(local_pes_19_16_io_out_sum),
    .io_out_sum_exp(local_pes_19_16_io_out_sum_exp),
    .io_out_kv(local_pes_19_16_io_out_kv),
    .io_out_stage(local_pes_19_16_io_out_stage)
  );
  PE_1 local_pes_19_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_17_clock),
    .reset(local_pes_19_17_reset),
    .io_in_q(local_pes_19_17_io_in_q),
    .io_in_sum(local_pes_19_17_io_in_sum),
    .io_in_sum_exp(local_pes_19_17_io_in_sum_exp),
    .io_in_kv(local_pes_19_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_17_io_in_inv_sum),
    .io_in_stage(local_pes_19_17_io_in_stage),
    .io_out_q(local_pes_19_17_io_out_q),
    .io_out_sum(local_pes_19_17_io_out_sum),
    .io_out_sum_exp(local_pes_19_17_io_out_sum_exp),
    .io_out_kv(local_pes_19_17_io_out_kv),
    .io_out_stage(local_pes_19_17_io_out_stage)
  );
  PE_1 local_pes_19_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_18_clock),
    .reset(local_pes_19_18_reset),
    .io_in_q(local_pes_19_18_io_in_q),
    .io_in_sum(local_pes_19_18_io_in_sum),
    .io_in_sum_exp(local_pes_19_18_io_in_sum_exp),
    .io_in_kv(local_pes_19_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_18_io_in_inv_sum),
    .io_in_stage(local_pes_19_18_io_in_stage),
    .io_out_q(local_pes_19_18_io_out_q),
    .io_out_sum(local_pes_19_18_io_out_sum),
    .io_out_sum_exp(local_pes_19_18_io_out_sum_exp),
    .io_out_kv(local_pes_19_18_io_out_kv),
    .io_out_stage(local_pes_19_18_io_out_stage)
  );
  PE_1 local_pes_19_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_19_clock),
    .reset(local_pes_19_19_reset),
    .io_in_q(local_pes_19_19_io_in_q),
    .io_in_sum(local_pes_19_19_io_in_sum),
    .io_in_sum_exp(local_pes_19_19_io_in_sum_exp),
    .io_in_kv(local_pes_19_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_19_io_in_inv_sum),
    .io_in_stage(local_pes_19_19_io_in_stage),
    .io_out_q(local_pes_19_19_io_out_q),
    .io_out_sum(local_pes_19_19_io_out_sum),
    .io_out_sum_exp(local_pes_19_19_io_out_sum_exp),
    .io_out_kv(local_pes_19_19_io_out_kv),
    .io_out_stage(local_pes_19_19_io_out_stage)
  );
  PE_1 local_pes_19_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_20_clock),
    .reset(local_pes_19_20_reset),
    .io_in_q(local_pes_19_20_io_in_q),
    .io_in_sum(local_pes_19_20_io_in_sum),
    .io_in_sum_exp(local_pes_19_20_io_in_sum_exp),
    .io_in_kv(local_pes_19_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_20_io_in_inv_sum),
    .io_in_stage(local_pes_19_20_io_in_stage),
    .io_out_q(local_pes_19_20_io_out_q),
    .io_out_sum(local_pes_19_20_io_out_sum),
    .io_out_sum_exp(local_pes_19_20_io_out_sum_exp),
    .io_out_kv(local_pes_19_20_io_out_kv),
    .io_out_stage(local_pes_19_20_io_out_stage)
  );
  PE_1 local_pes_19_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_21_clock),
    .reset(local_pes_19_21_reset),
    .io_in_q(local_pes_19_21_io_in_q),
    .io_in_sum(local_pes_19_21_io_in_sum),
    .io_in_sum_exp(local_pes_19_21_io_in_sum_exp),
    .io_in_kv(local_pes_19_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_21_io_in_inv_sum),
    .io_in_stage(local_pes_19_21_io_in_stage),
    .io_out_q(local_pes_19_21_io_out_q),
    .io_out_sum(local_pes_19_21_io_out_sum),
    .io_out_sum_exp(local_pes_19_21_io_out_sum_exp),
    .io_out_kv(local_pes_19_21_io_out_kv),
    .io_out_stage(local_pes_19_21_io_out_stage)
  );
  PE_1 local_pes_19_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_22_clock),
    .reset(local_pes_19_22_reset),
    .io_in_q(local_pes_19_22_io_in_q),
    .io_in_sum(local_pes_19_22_io_in_sum),
    .io_in_sum_exp(local_pes_19_22_io_in_sum_exp),
    .io_in_kv(local_pes_19_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_22_io_in_inv_sum),
    .io_in_stage(local_pes_19_22_io_in_stage),
    .io_out_q(local_pes_19_22_io_out_q),
    .io_out_sum(local_pes_19_22_io_out_sum),
    .io_out_sum_exp(local_pes_19_22_io_out_sum_exp),
    .io_out_kv(local_pes_19_22_io_out_kv),
    .io_out_stage(local_pes_19_22_io_out_stage)
  );
  PE_1 local_pes_19_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_23_clock),
    .reset(local_pes_19_23_reset),
    .io_in_q(local_pes_19_23_io_in_q),
    .io_in_sum(local_pes_19_23_io_in_sum),
    .io_in_sum_exp(local_pes_19_23_io_in_sum_exp),
    .io_in_kv(local_pes_19_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_23_io_in_inv_sum),
    .io_in_stage(local_pes_19_23_io_in_stage),
    .io_out_q(local_pes_19_23_io_out_q),
    .io_out_sum(local_pes_19_23_io_out_sum),
    .io_out_sum_exp(local_pes_19_23_io_out_sum_exp),
    .io_out_kv(local_pes_19_23_io_out_kv),
    .io_out_stage(local_pes_19_23_io_out_stage)
  );
  PE_1 local_pes_19_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_24_clock),
    .reset(local_pes_19_24_reset),
    .io_in_q(local_pes_19_24_io_in_q),
    .io_in_sum(local_pes_19_24_io_in_sum),
    .io_in_sum_exp(local_pes_19_24_io_in_sum_exp),
    .io_in_kv(local_pes_19_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_24_io_in_inv_sum),
    .io_in_stage(local_pes_19_24_io_in_stage),
    .io_out_q(local_pes_19_24_io_out_q),
    .io_out_sum(local_pes_19_24_io_out_sum),
    .io_out_sum_exp(local_pes_19_24_io_out_sum_exp),
    .io_out_kv(local_pes_19_24_io_out_kv),
    .io_out_stage(local_pes_19_24_io_out_stage)
  );
  PE_1 local_pes_19_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_25_clock),
    .reset(local_pes_19_25_reset),
    .io_in_q(local_pes_19_25_io_in_q),
    .io_in_sum(local_pes_19_25_io_in_sum),
    .io_in_sum_exp(local_pes_19_25_io_in_sum_exp),
    .io_in_kv(local_pes_19_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_25_io_in_inv_sum),
    .io_in_stage(local_pes_19_25_io_in_stage),
    .io_out_q(local_pes_19_25_io_out_q),
    .io_out_sum(local_pes_19_25_io_out_sum),
    .io_out_sum_exp(local_pes_19_25_io_out_sum_exp),
    .io_out_kv(local_pes_19_25_io_out_kv),
    .io_out_stage(local_pes_19_25_io_out_stage)
  );
  PE_1 local_pes_19_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_26_clock),
    .reset(local_pes_19_26_reset),
    .io_in_q(local_pes_19_26_io_in_q),
    .io_in_sum(local_pes_19_26_io_in_sum),
    .io_in_sum_exp(local_pes_19_26_io_in_sum_exp),
    .io_in_kv(local_pes_19_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_26_io_in_inv_sum),
    .io_in_stage(local_pes_19_26_io_in_stage),
    .io_out_q(local_pes_19_26_io_out_q),
    .io_out_sum(local_pes_19_26_io_out_sum),
    .io_out_sum_exp(local_pes_19_26_io_out_sum_exp),
    .io_out_kv(local_pes_19_26_io_out_kv),
    .io_out_stage(local_pes_19_26_io_out_stage)
  );
  PE_1 local_pes_19_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_27_clock),
    .reset(local_pes_19_27_reset),
    .io_in_q(local_pes_19_27_io_in_q),
    .io_in_sum(local_pes_19_27_io_in_sum),
    .io_in_sum_exp(local_pes_19_27_io_in_sum_exp),
    .io_in_kv(local_pes_19_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_27_io_in_inv_sum),
    .io_in_stage(local_pes_19_27_io_in_stage),
    .io_out_q(local_pes_19_27_io_out_q),
    .io_out_sum(local_pes_19_27_io_out_sum),
    .io_out_sum_exp(local_pes_19_27_io_out_sum_exp),
    .io_out_kv(local_pes_19_27_io_out_kv),
    .io_out_stage(local_pes_19_27_io_out_stage)
  );
  PE_1 local_pes_19_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_28_clock),
    .reset(local_pes_19_28_reset),
    .io_in_q(local_pes_19_28_io_in_q),
    .io_in_sum(local_pes_19_28_io_in_sum),
    .io_in_sum_exp(local_pes_19_28_io_in_sum_exp),
    .io_in_kv(local_pes_19_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_28_io_in_inv_sum),
    .io_in_stage(local_pes_19_28_io_in_stage),
    .io_out_q(local_pes_19_28_io_out_q),
    .io_out_sum(local_pes_19_28_io_out_sum),
    .io_out_sum_exp(local_pes_19_28_io_out_sum_exp),
    .io_out_kv(local_pes_19_28_io_out_kv),
    .io_out_stage(local_pes_19_28_io_out_stage)
  );
  PE_1 local_pes_19_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_29_clock),
    .reset(local_pes_19_29_reset),
    .io_in_q(local_pes_19_29_io_in_q),
    .io_in_sum(local_pes_19_29_io_in_sum),
    .io_in_sum_exp(local_pes_19_29_io_in_sum_exp),
    .io_in_kv(local_pes_19_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_29_io_in_inv_sum),
    .io_in_stage(local_pes_19_29_io_in_stage),
    .io_out_q(local_pes_19_29_io_out_q),
    .io_out_sum(local_pes_19_29_io_out_sum),
    .io_out_sum_exp(local_pes_19_29_io_out_sum_exp),
    .io_out_kv(local_pes_19_29_io_out_kv),
    .io_out_stage(local_pes_19_29_io_out_stage)
  );
  PE_1 local_pes_19_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_30_clock),
    .reset(local_pes_19_30_reset),
    .io_in_q(local_pes_19_30_io_in_q),
    .io_in_sum(local_pes_19_30_io_in_sum),
    .io_in_sum_exp(local_pes_19_30_io_in_sum_exp),
    .io_in_kv(local_pes_19_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_30_io_in_inv_sum),
    .io_in_stage(local_pes_19_30_io_in_stage),
    .io_out_q(local_pes_19_30_io_out_q),
    .io_out_sum(local_pes_19_30_io_out_sum),
    .io_out_sum_exp(local_pes_19_30_io_out_sum_exp),
    .io_out_kv(local_pes_19_30_io_out_kv),
    .io_out_stage(local_pes_19_30_io_out_stage)
  );
  PE_1 local_pes_19_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_19_31_clock),
    .reset(local_pes_19_31_reset),
    .io_in_q(local_pes_19_31_io_in_q),
    .io_in_sum(local_pes_19_31_io_in_sum),
    .io_in_sum_exp(local_pes_19_31_io_in_sum_exp),
    .io_in_kv(local_pes_19_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_19_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_19_31_io_in_inv_sum),
    .io_in_stage(local_pes_19_31_io_in_stage),
    .io_out_q(local_pes_19_31_io_out_q),
    .io_out_sum(local_pes_19_31_io_out_sum),
    .io_out_sum_exp(local_pes_19_31_io_out_sum_exp),
    .io_out_kv(local_pes_19_31_io_out_kv),
    .io_out_stage(local_pes_19_31_io_out_stage)
  );
  PE local_pes_20_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_0_clock),
    .reset(local_pes_20_0_reset),
    .io_in_q(local_pes_20_0_io_in_q),
    .io_in_kv(local_pes_20_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_0_io_in_inv_sum),
    .io_in_stage(local_pes_20_0_io_in_stage),
    .io_out_q(local_pes_20_0_io_out_q),
    .io_out_sum(local_pes_20_0_io_out_sum),
    .io_out_kv(local_pes_20_0_io_out_kv),
    .io_out_stage(local_pes_20_0_io_out_stage)
  );
  PE_1 local_pes_20_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_1_clock),
    .reset(local_pes_20_1_reset),
    .io_in_q(local_pes_20_1_io_in_q),
    .io_in_sum(local_pes_20_1_io_in_sum),
    .io_in_sum_exp(local_pes_20_1_io_in_sum_exp),
    .io_in_kv(local_pes_20_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_1_io_in_inv_sum),
    .io_in_stage(local_pes_20_1_io_in_stage),
    .io_out_q(local_pes_20_1_io_out_q),
    .io_out_sum(local_pes_20_1_io_out_sum),
    .io_out_sum_exp(local_pes_20_1_io_out_sum_exp),
    .io_out_kv(local_pes_20_1_io_out_kv),
    .io_out_stage(local_pes_20_1_io_out_stage)
  );
  PE_1 local_pes_20_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_2_clock),
    .reset(local_pes_20_2_reset),
    .io_in_q(local_pes_20_2_io_in_q),
    .io_in_sum(local_pes_20_2_io_in_sum),
    .io_in_sum_exp(local_pes_20_2_io_in_sum_exp),
    .io_in_kv(local_pes_20_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_2_io_in_inv_sum),
    .io_in_stage(local_pes_20_2_io_in_stage),
    .io_out_q(local_pes_20_2_io_out_q),
    .io_out_sum(local_pes_20_2_io_out_sum),
    .io_out_sum_exp(local_pes_20_2_io_out_sum_exp),
    .io_out_kv(local_pes_20_2_io_out_kv),
    .io_out_stage(local_pes_20_2_io_out_stage)
  );
  PE_1 local_pes_20_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_3_clock),
    .reset(local_pes_20_3_reset),
    .io_in_q(local_pes_20_3_io_in_q),
    .io_in_sum(local_pes_20_3_io_in_sum),
    .io_in_sum_exp(local_pes_20_3_io_in_sum_exp),
    .io_in_kv(local_pes_20_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_3_io_in_inv_sum),
    .io_in_stage(local_pes_20_3_io_in_stage),
    .io_out_q(local_pes_20_3_io_out_q),
    .io_out_sum(local_pes_20_3_io_out_sum),
    .io_out_sum_exp(local_pes_20_3_io_out_sum_exp),
    .io_out_kv(local_pes_20_3_io_out_kv),
    .io_out_stage(local_pes_20_3_io_out_stage)
  );
  PE_1 local_pes_20_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_4_clock),
    .reset(local_pes_20_4_reset),
    .io_in_q(local_pes_20_4_io_in_q),
    .io_in_sum(local_pes_20_4_io_in_sum),
    .io_in_sum_exp(local_pes_20_4_io_in_sum_exp),
    .io_in_kv(local_pes_20_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_4_io_in_inv_sum),
    .io_in_stage(local_pes_20_4_io_in_stage),
    .io_out_q(local_pes_20_4_io_out_q),
    .io_out_sum(local_pes_20_4_io_out_sum),
    .io_out_sum_exp(local_pes_20_4_io_out_sum_exp),
    .io_out_kv(local_pes_20_4_io_out_kv),
    .io_out_stage(local_pes_20_4_io_out_stage)
  );
  PE_1 local_pes_20_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_5_clock),
    .reset(local_pes_20_5_reset),
    .io_in_q(local_pes_20_5_io_in_q),
    .io_in_sum(local_pes_20_5_io_in_sum),
    .io_in_sum_exp(local_pes_20_5_io_in_sum_exp),
    .io_in_kv(local_pes_20_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_5_io_in_inv_sum),
    .io_in_stage(local_pes_20_5_io_in_stage),
    .io_out_q(local_pes_20_5_io_out_q),
    .io_out_sum(local_pes_20_5_io_out_sum),
    .io_out_sum_exp(local_pes_20_5_io_out_sum_exp),
    .io_out_kv(local_pes_20_5_io_out_kv),
    .io_out_stage(local_pes_20_5_io_out_stage)
  );
  PE_1 local_pes_20_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_6_clock),
    .reset(local_pes_20_6_reset),
    .io_in_q(local_pes_20_6_io_in_q),
    .io_in_sum(local_pes_20_6_io_in_sum),
    .io_in_sum_exp(local_pes_20_6_io_in_sum_exp),
    .io_in_kv(local_pes_20_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_6_io_in_inv_sum),
    .io_in_stage(local_pes_20_6_io_in_stage),
    .io_out_q(local_pes_20_6_io_out_q),
    .io_out_sum(local_pes_20_6_io_out_sum),
    .io_out_sum_exp(local_pes_20_6_io_out_sum_exp),
    .io_out_kv(local_pes_20_6_io_out_kv),
    .io_out_stage(local_pes_20_6_io_out_stage)
  );
  PE_1 local_pes_20_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_7_clock),
    .reset(local_pes_20_7_reset),
    .io_in_q(local_pes_20_7_io_in_q),
    .io_in_sum(local_pes_20_7_io_in_sum),
    .io_in_sum_exp(local_pes_20_7_io_in_sum_exp),
    .io_in_kv(local_pes_20_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_7_io_in_inv_sum),
    .io_in_stage(local_pes_20_7_io_in_stage),
    .io_out_q(local_pes_20_7_io_out_q),
    .io_out_sum(local_pes_20_7_io_out_sum),
    .io_out_sum_exp(local_pes_20_7_io_out_sum_exp),
    .io_out_kv(local_pes_20_7_io_out_kv),
    .io_out_stage(local_pes_20_7_io_out_stage)
  );
  PE_1 local_pes_20_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_8_clock),
    .reset(local_pes_20_8_reset),
    .io_in_q(local_pes_20_8_io_in_q),
    .io_in_sum(local_pes_20_8_io_in_sum),
    .io_in_sum_exp(local_pes_20_8_io_in_sum_exp),
    .io_in_kv(local_pes_20_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_8_io_in_inv_sum),
    .io_in_stage(local_pes_20_8_io_in_stage),
    .io_out_q(local_pes_20_8_io_out_q),
    .io_out_sum(local_pes_20_8_io_out_sum),
    .io_out_sum_exp(local_pes_20_8_io_out_sum_exp),
    .io_out_kv(local_pes_20_8_io_out_kv),
    .io_out_stage(local_pes_20_8_io_out_stage)
  );
  PE_1 local_pes_20_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_9_clock),
    .reset(local_pes_20_9_reset),
    .io_in_q(local_pes_20_9_io_in_q),
    .io_in_sum(local_pes_20_9_io_in_sum),
    .io_in_sum_exp(local_pes_20_9_io_in_sum_exp),
    .io_in_kv(local_pes_20_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_9_io_in_inv_sum),
    .io_in_stage(local_pes_20_9_io_in_stage),
    .io_out_q(local_pes_20_9_io_out_q),
    .io_out_sum(local_pes_20_9_io_out_sum),
    .io_out_sum_exp(local_pes_20_9_io_out_sum_exp),
    .io_out_kv(local_pes_20_9_io_out_kv),
    .io_out_stage(local_pes_20_9_io_out_stage)
  );
  PE_1 local_pes_20_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_10_clock),
    .reset(local_pes_20_10_reset),
    .io_in_q(local_pes_20_10_io_in_q),
    .io_in_sum(local_pes_20_10_io_in_sum),
    .io_in_sum_exp(local_pes_20_10_io_in_sum_exp),
    .io_in_kv(local_pes_20_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_10_io_in_inv_sum),
    .io_in_stage(local_pes_20_10_io_in_stage),
    .io_out_q(local_pes_20_10_io_out_q),
    .io_out_sum(local_pes_20_10_io_out_sum),
    .io_out_sum_exp(local_pes_20_10_io_out_sum_exp),
    .io_out_kv(local_pes_20_10_io_out_kv),
    .io_out_stage(local_pes_20_10_io_out_stage)
  );
  PE_1 local_pes_20_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_11_clock),
    .reset(local_pes_20_11_reset),
    .io_in_q(local_pes_20_11_io_in_q),
    .io_in_sum(local_pes_20_11_io_in_sum),
    .io_in_sum_exp(local_pes_20_11_io_in_sum_exp),
    .io_in_kv(local_pes_20_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_11_io_in_inv_sum),
    .io_in_stage(local_pes_20_11_io_in_stage),
    .io_out_q(local_pes_20_11_io_out_q),
    .io_out_sum(local_pes_20_11_io_out_sum),
    .io_out_sum_exp(local_pes_20_11_io_out_sum_exp),
    .io_out_kv(local_pes_20_11_io_out_kv),
    .io_out_stage(local_pes_20_11_io_out_stage)
  );
  PE_1 local_pes_20_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_12_clock),
    .reset(local_pes_20_12_reset),
    .io_in_q(local_pes_20_12_io_in_q),
    .io_in_sum(local_pes_20_12_io_in_sum),
    .io_in_sum_exp(local_pes_20_12_io_in_sum_exp),
    .io_in_kv(local_pes_20_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_12_io_in_inv_sum),
    .io_in_stage(local_pes_20_12_io_in_stage),
    .io_out_q(local_pes_20_12_io_out_q),
    .io_out_sum(local_pes_20_12_io_out_sum),
    .io_out_sum_exp(local_pes_20_12_io_out_sum_exp),
    .io_out_kv(local_pes_20_12_io_out_kv),
    .io_out_stage(local_pes_20_12_io_out_stage)
  );
  PE_1 local_pes_20_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_13_clock),
    .reset(local_pes_20_13_reset),
    .io_in_q(local_pes_20_13_io_in_q),
    .io_in_sum(local_pes_20_13_io_in_sum),
    .io_in_sum_exp(local_pes_20_13_io_in_sum_exp),
    .io_in_kv(local_pes_20_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_13_io_in_inv_sum),
    .io_in_stage(local_pes_20_13_io_in_stage),
    .io_out_q(local_pes_20_13_io_out_q),
    .io_out_sum(local_pes_20_13_io_out_sum),
    .io_out_sum_exp(local_pes_20_13_io_out_sum_exp),
    .io_out_kv(local_pes_20_13_io_out_kv),
    .io_out_stage(local_pes_20_13_io_out_stage)
  );
  PE_1 local_pes_20_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_14_clock),
    .reset(local_pes_20_14_reset),
    .io_in_q(local_pes_20_14_io_in_q),
    .io_in_sum(local_pes_20_14_io_in_sum),
    .io_in_sum_exp(local_pes_20_14_io_in_sum_exp),
    .io_in_kv(local_pes_20_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_14_io_in_inv_sum),
    .io_in_stage(local_pes_20_14_io_in_stage),
    .io_out_q(local_pes_20_14_io_out_q),
    .io_out_sum(local_pes_20_14_io_out_sum),
    .io_out_sum_exp(local_pes_20_14_io_out_sum_exp),
    .io_out_kv(local_pes_20_14_io_out_kv),
    .io_out_stage(local_pes_20_14_io_out_stage)
  );
  PE_1 local_pes_20_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_15_clock),
    .reset(local_pes_20_15_reset),
    .io_in_q(local_pes_20_15_io_in_q),
    .io_in_sum(local_pes_20_15_io_in_sum),
    .io_in_sum_exp(local_pes_20_15_io_in_sum_exp),
    .io_in_kv(local_pes_20_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_15_io_in_inv_sum),
    .io_in_stage(local_pes_20_15_io_in_stage),
    .io_out_q(local_pes_20_15_io_out_q),
    .io_out_sum(local_pes_20_15_io_out_sum),
    .io_out_sum_exp(local_pes_20_15_io_out_sum_exp),
    .io_out_kv(local_pes_20_15_io_out_kv),
    .io_out_stage(local_pes_20_15_io_out_stage)
  );
  PE_1 local_pes_20_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_16_clock),
    .reset(local_pes_20_16_reset),
    .io_in_q(local_pes_20_16_io_in_q),
    .io_in_sum(local_pes_20_16_io_in_sum),
    .io_in_sum_exp(local_pes_20_16_io_in_sum_exp),
    .io_in_kv(local_pes_20_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_16_io_in_inv_sum),
    .io_in_stage(local_pes_20_16_io_in_stage),
    .io_out_q(local_pes_20_16_io_out_q),
    .io_out_sum(local_pes_20_16_io_out_sum),
    .io_out_sum_exp(local_pes_20_16_io_out_sum_exp),
    .io_out_kv(local_pes_20_16_io_out_kv),
    .io_out_stage(local_pes_20_16_io_out_stage)
  );
  PE_1 local_pes_20_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_17_clock),
    .reset(local_pes_20_17_reset),
    .io_in_q(local_pes_20_17_io_in_q),
    .io_in_sum(local_pes_20_17_io_in_sum),
    .io_in_sum_exp(local_pes_20_17_io_in_sum_exp),
    .io_in_kv(local_pes_20_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_17_io_in_inv_sum),
    .io_in_stage(local_pes_20_17_io_in_stage),
    .io_out_q(local_pes_20_17_io_out_q),
    .io_out_sum(local_pes_20_17_io_out_sum),
    .io_out_sum_exp(local_pes_20_17_io_out_sum_exp),
    .io_out_kv(local_pes_20_17_io_out_kv),
    .io_out_stage(local_pes_20_17_io_out_stage)
  );
  PE_1 local_pes_20_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_18_clock),
    .reset(local_pes_20_18_reset),
    .io_in_q(local_pes_20_18_io_in_q),
    .io_in_sum(local_pes_20_18_io_in_sum),
    .io_in_sum_exp(local_pes_20_18_io_in_sum_exp),
    .io_in_kv(local_pes_20_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_18_io_in_inv_sum),
    .io_in_stage(local_pes_20_18_io_in_stage),
    .io_out_q(local_pes_20_18_io_out_q),
    .io_out_sum(local_pes_20_18_io_out_sum),
    .io_out_sum_exp(local_pes_20_18_io_out_sum_exp),
    .io_out_kv(local_pes_20_18_io_out_kv),
    .io_out_stage(local_pes_20_18_io_out_stage)
  );
  PE_1 local_pes_20_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_19_clock),
    .reset(local_pes_20_19_reset),
    .io_in_q(local_pes_20_19_io_in_q),
    .io_in_sum(local_pes_20_19_io_in_sum),
    .io_in_sum_exp(local_pes_20_19_io_in_sum_exp),
    .io_in_kv(local_pes_20_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_19_io_in_inv_sum),
    .io_in_stage(local_pes_20_19_io_in_stage),
    .io_out_q(local_pes_20_19_io_out_q),
    .io_out_sum(local_pes_20_19_io_out_sum),
    .io_out_sum_exp(local_pes_20_19_io_out_sum_exp),
    .io_out_kv(local_pes_20_19_io_out_kv),
    .io_out_stage(local_pes_20_19_io_out_stage)
  );
  PE_1 local_pes_20_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_20_clock),
    .reset(local_pes_20_20_reset),
    .io_in_q(local_pes_20_20_io_in_q),
    .io_in_sum(local_pes_20_20_io_in_sum),
    .io_in_sum_exp(local_pes_20_20_io_in_sum_exp),
    .io_in_kv(local_pes_20_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_20_io_in_inv_sum),
    .io_in_stage(local_pes_20_20_io_in_stage),
    .io_out_q(local_pes_20_20_io_out_q),
    .io_out_sum(local_pes_20_20_io_out_sum),
    .io_out_sum_exp(local_pes_20_20_io_out_sum_exp),
    .io_out_kv(local_pes_20_20_io_out_kv),
    .io_out_stage(local_pes_20_20_io_out_stage)
  );
  PE_1 local_pes_20_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_21_clock),
    .reset(local_pes_20_21_reset),
    .io_in_q(local_pes_20_21_io_in_q),
    .io_in_sum(local_pes_20_21_io_in_sum),
    .io_in_sum_exp(local_pes_20_21_io_in_sum_exp),
    .io_in_kv(local_pes_20_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_21_io_in_inv_sum),
    .io_in_stage(local_pes_20_21_io_in_stage),
    .io_out_q(local_pes_20_21_io_out_q),
    .io_out_sum(local_pes_20_21_io_out_sum),
    .io_out_sum_exp(local_pes_20_21_io_out_sum_exp),
    .io_out_kv(local_pes_20_21_io_out_kv),
    .io_out_stage(local_pes_20_21_io_out_stage)
  );
  PE_1 local_pes_20_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_22_clock),
    .reset(local_pes_20_22_reset),
    .io_in_q(local_pes_20_22_io_in_q),
    .io_in_sum(local_pes_20_22_io_in_sum),
    .io_in_sum_exp(local_pes_20_22_io_in_sum_exp),
    .io_in_kv(local_pes_20_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_22_io_in_inv_sum),
    .io_in_stage(local_pes_20_22_io_in_stage),
    .io_out_q(local_pes_20_22_io_out_q),
    .io_out_sum(local_pes_20_22_io_out_sum),
    .io_out_sum_exp(local_pes_20_22_io_out_sum_exp),
    .io_out_kv(local_pes_20_22_io_out_kv),
    .io_out_stage(local_pes_20_22_io_out_stage)
  );
  PE_1 local_pes_20_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_23_clock),
    .reset(local_pes_20_23_reset),
    .io_in_q(local_pes_20_23_io_in_q),
    .io_in_sum(local_pes_20_23_io_in_sum),
    .io_in_sum_exp(local_pes_20_23_io_in_sum_exp),
    .io_in_kv(local_pes_20_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_23_io_in_inv_sum),
    .io_in_stage(local_pes_20_23_io_in_stage),
    .io_out_q(local_pes_20_23_io_out_q),
    .io_out_sum(local_pes_20_23_io_out_sum),
    .io_out_sum_exp(local_pes_20_23_io_out_sum_exp),
    .io_out_kv(local_pes_20_23_io_out_kv),
    .io_out_stage(local_pes_20_23_io_out_stage)
  );
  PE_1 local_pes_20_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_24_clock),
    .reset(local_pes_20_24_reset),
    .io_in_q(local_pes_20_24_io_in_q),
    .io_in_sum(local_pes_20_24_io_in_sum),
    .io_in_sum_exp(local_pes_20_24_io_in_sum_exp),
    .io_in_kv(local_pes_20_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_24_io_in_inv_sum),
    .io_in_stage(local_pes_20_24_io_in_stage),
    .io_out_q(local_pes_20_24_io_out_q),
    .io_out_sum(local_pes_20_24_io_out_sum),
    .io_out_sum_exp(local_pes_20_24_io_out_sum_exp),
    .io_out_kv(local_pes_20_24_io_out_kv),
    .io_out_stage(local_pes_20_24_io_out_stage)
  );
  PE_1 local_pes_20_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_25_clock),
    .reset(local_pes_20_25_reset),
    .io_in_q(local_pes_20_25_io_in_q),
    .io_in_sum(local_pes_20_25_io_in_sum),
    .io_in_sum_exp(local_pes_20_25_io_in_sum_exp),
    .io_in_kv(local_pes_20_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_25_io_in_inv_sum),
    .io_in_stage(local_pes_20_25_io_in_stage),
    .io_out_q(local_pes_20_25_io_out_q),
    .io_out_sum(local_pes_20_25_io_out_sum),
    .io_out_sum_exp(local_pes_20_25_io_out_sum_exp),
    .io_out_kv(local_pes_20_25_io_out_kv),
    .io_out_stage(local_pes_20_25_io_out_stage)
  );
  PE_1 local_pes_20_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_26_clock),
    .reset(local_pes_20_26_reset),
    .io_in_q(local_pes_20_26_io_in_q),
    .io_in_sum(local_pes_20_26_io_in_sum),
    .io_in_sum_exp(local_pes_20_26_io_in_sum_exp),
    .io_in_kv(local_pes_20_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_26_io_in_inv_sum),
    .io_in_stage(local_pes_20_26_io_in_stage),
    .io_out_q(local_pes_20_26_io_out_q),
    .io_out_sum(local_pes_20_26_io_out_sum),
    .io_out_sum_exp(local_pes_20_26_io_out_sum_exp),
    .io_out_kv(local_pes_20_26_io_out_kv),
    .io_out_stage(local_pes_20_26_io_out_stage)
  );
  PE_1 local_pes_20_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_27_clock),
    .reset(local_pes_20_27_reset),
    .io_in_q(local_pes_20_27_io_in_q),
    .io_in_sum(local_pes_20_27_io_in_sum),
    .io_in_sum_exp(local_pes_20_27_io_in_sum_exp),
    .io_in_kv(local_pes_20_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_27_io_in_inv_sum),
    .io_in_stage(local_pes_20_27_io_in_stage),
    .io_out_q(local_pes_20_27_io_out_q),
    .io_out_sum(local_pes_20_27_io_out_sum),
    .io_out_sum_exp(local_pes_20_27_io_out_sum_exp),
    .io_out_kv(local_pes_20_27_io_out_kv),
    .io_out_stage(local_pes_20_27_io_out_stage)
  );
  PE_1 local_pes_20_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_28_clock),
    .reset(local_pes_20_28_reset),
    .io_in_q(local_pes_20_28_io_in_q),
    .io_in_sum(local_pes_20_28_io_in_sum),
    .io_in_sum_exp(local_pes_20_28_io_in_sum_exp),
    .io_in_kv(local_pes_20_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_28_io_in_inv_sum),
    .io_in_stage(local_pes_20_28_io_in_stage),
    .io_out_q(local_pes_20_28_io_out_q),
    .io_out_sum(local_pes_20_28_io_out_sum),
    .io_out_sum_exp(local_pes_20_28_io_out_sum_exp),
    .io_out_kv(local_pes_20_28_io_out_kv),
    .io_out_stage(local_pes_20_28_io_out_stage)
  );
  PE_1 local_pes_20_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_29_clock),
    .reset(local_pes_20_29_reset),
    .io_in_q(local_pes_20_29_io_in_q),
    .io_in_sum(local_pes_20_29_io_in_sum),
    .io_in_sum_exp(local_pes_20_29_io_in_sum_exp),
    .io_in_kv(local_pes_20_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_29_io_in_inv_sum),
    .io_in_stage(local_pes_20_29_io_in_stage),
    .io_out_q(local_pes_20_29_io_out_q),
    .io_out_sum(local_pes_20_29_io_out_sum),
    .io_out_sum_exp(local_pes_20_29_io_out_sum_exp),
    .io_out_kv(local_pes_20_29_io_out_kv),
    .io_out_stage(local_pes_20_29_io_out_stage)
  );
  PE_1 local_pes_20_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_30_clock),
    .reset(local_pes_20_30_reset),
    .io_in_q(local_pes_20_30_io_in_q),
    .io_in_sum(local_pes_20_30_io_in_sum),
    .io_in_sum_exp(local_pes_20_30_io_in_sum_exp),
    .io_in_kv(local_pes_20_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_30_io_in_inv_sum),
    .io_in_stage(local_pes_20_30_io_in_stage),
    .io_out_q(local_pes_20_30_io_out_q),
    .io_out_sum(local_pes_20_30_io_out_sum),
    .io_out_sum_exp(local_pes_20_30_io_out_sum_exp),
    .io_out_kv(local_pes_20_30_io_out_kv),
    .io_out_stage(local_pes_20_30_io_out_stage)
  );
  PE_1 local_pes_20_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_20_31_clock),
    .reset(local_pes_20_31_reset),
    .io_in_q(local_pes_20_31_io_in_q),
    .io_in_sum(local_pes_20_31_io_in_sum),
    .io_in_sum_exp(local_pes_20_31_io_in_sum_exp),
    .io_in_kv(local_pes_20_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_20_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_20_31_io_in_inv_sum),
    .io_in_stage(local_pes_20_31_io_in_stage),
    .io_out_q(local_pes_20_31_io_out_q),
    .io_out_sum(local_pes_20_31_io_out_sum),
    .io_out_sum_exp(local_pes_20_31_io_out_sum_exp),
    .io_out_kv(local_pes_20_31_io_out_kv),
    .io_out_stage(local_pes_20_31_io_out_stage)
  );
  PE local_pes_21_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_0_clock),
    .reset(local_pes_21_0_reset),
    .io_in_q(local_pes_21_0_io_in_q),
    .io_in_kv(local_pes_21_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_0_io_in_inv_sum),
    .io_in_stage(local_pes_21_0_io_in_stage),
    .io_out_q(local_pes_21_0_io_out_q),
    .io_out_sum(local_pes_21_0_io_out_sum),
    .io_out_kv(local_pes_21_0_io_out_kv),
    .io_out_stage(local_pes_21_0_io_out_stage)
  );
  PE_1 local_pes_21_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_1_clock),
    .reset(local_pes_21_1_reset),
    .io_in_q(local_pes_21_1_io_in_q),
    .io_in_sum(local_pes_21_1_io_in_sum),
    .io_in_sum_exp(local_pes_21_1_io_in_sum_exp),
    .io_in_kv(local_pes_21_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_1_io_in_inv_sum),
    .io_in_stage(local_pes_21_1_io_in_stage),
    .io_out_q(local_pes_21_1_io_out_q),
    .io_out_sum(local_pes_21_1_io_out_sum),
    .io_out_sum_exp(local_pes_21_1_io_out_sum_exp),
    .io_out_kv(local_pes_21_1_io_out_kv),
    .io_out_stage(local_pes_21_1_io_out_stage)
  );
  PE_1 local_pes_21_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_2_clock),
    .reset(local_pes_21_2_reset),
    .io_in_q(local_pes_21_2_io_in_q),
    .io_in_sum(local_pes_21_2_io_in_sum),
    .io_in_sum_exp(local_pes_21_2_io_in_sum_exp),
    .io_in_kv(local_pes_21_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_2_io_in_inv_sum),
    .io_in_stage(local_pes_21_2_io_in_stage),
    .io_out_q(local_pes_21_2_io_out_q),
    .io_out_sum(local_pes_21_2_io_out_sum),
    .io_out_sum_exp(local_pes_21_2_io_out_sum_exp),
    .io_out_kv(local_pes_21_2_io_out_kv),
    .io_out_stage(local_pes_21_2_io_out_stage)
  );
  PE_1 local_pes_21_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_3_clock),
    .reset(local_pes_21_3_reset),
    .io_in_q(local_pes_21_3_io_in_q),
    .io_in_sum(local_pes_21_3_io_in_sum),
    .io_in_sum_exp(local_pes_21_3_io_in_sum_exp),
    .io_in_kv(local_pes_21_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_3_io_in_inv_sum),
    .io_in_stage(local_pes_21_3_io_in_stage),
    .io_out_q(local_pes_21_3_io_out_q),
    .io_out_sum(local_pes_21_3_io_out_sum),
    .io_out_sum_exp(local_pes_21_3_io_out_sum_exp),
    .io_out_kv(local_pes_21_3_io_out_kv),
    .io_out_stage(local_pes_21_3_io_out_stage)
  );
  PE_1 local_pes_21_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_4_clock),
    .reset(local_pes_21_4_reset),
    .io_in_q(local_pes_21_4_io_in_q),
    .io_in_sum(local_pes_21_4_io_in_sum),
    .io_in_sum_exp(local_pes_21_4_io_in_sum_exp),
    .io_in_kv(local_pes_21_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_4_io_in_inv_sum),
    .io_in_stage(local_pes_21_4_io_in_stage),
    .io_out_q(local_pes_21_4_io_out_q),
    .io_out_sum(local_pes_21_4_io_out_sum),
    .io_out_sum_exp(local_pes_21_4_io_out_sum_exp),
    .io_out_kv(local_pes_21_4_io_out_kv),
    .io_out_stage(local_pes_21_4_io_out_stage)
  );
  PE_1 local_pes_21_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_5_clock),
    .reset(local_pes_21_5_reset),
    .io_in_q(local_pes_21_5_io_in_q),
    .io_in_sum(local_pes_21_5_io_in_sum),
    .io_in_sum_exp(local_pes_21_5_io_in_sum_exp),
    .io_in_kv(local_pes_21_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_5_io_in_inv_sum),
    .io_in_stage(local_pes_21_5_io_in_stage),
    .io_out_q(local_pes_21_5_io_out_q),
    .io_out_sum(local_pes_21_5_io_out_sum),
    .io_out_sum_exp(local_pes_21_5_io_out_sum_exp),
    .io_out_kv(local_pes_21_5_io_out_kv),
    .io_out_stage(local_pes_21_5_io_out_stage)
  );
  PE_1 local_pes_21_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_6_clock),
    .reset(local_pes_21_6_reset),
    .io_in_q(local_pes_21_6_io_in_q),
    .io_in_sum(local_pes_21_6_io_in_sum),
    .io_in_sum_exp(local_pes_21_6_io_in_sum_exp),
    .io_in_kv(local_pes_21_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_6_io_in_inv_sum),
    .io_in_stage(local_pes_21_6_io_in_stage),
    .io_out_q(local_pes_21_6_io_out_q),
    .io_out_sum(local_pes_21_6_io_out_sum),
    .io_out_sum_exp(local_pes_21_6_io_out_sum_exp),
    .io_out_kv(local_pes_21_6_io_out_kv),
    .io_out_stage(local_pes_21_6_io_out_stage)
  );
  PE_1 local_pes_21_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_7_clock),
    .reset(local_pes_21_7_reset),
    .io_in_q(local_pes_21_7_io_in_q),
    .io_in_sum(local_pes_21_7_io_in_sum),
    .io_in_sum_exp(local_pes_21_7_io_in_sum_exp),
    .io_in_kv(local_pes_21_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_7_io_in_inv_sum),
    .io_in_stage(local_pes_21_7_io_in_stage),
    .io_out_q(local_pes_21_7_io_out_q),
    .io_out_sum(local_pes_21_7_io_out_sum),
    .io_out_sum_exp(local_pes_21_7_io_out_sum_exp),
    .io_out_kv(local_pes_21_7_io_out_kv),
    .io_out_stage(local_pes_21_7_io_out_stage)
  );
  PE_1 local_pes_21_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_8_clock),
    .reset(local_pes_21_8_reset),
    .io_in_q(local_pes_21_8_io_in_q),
    .io_in_sum(local_pes_21_8_io_in_sum),
    .io_in_sum_exp(local_pes_21_8_io_in_sum_exp),
    .io_in_kv(local_pes_21_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_8_io_in_inv_sum),
    .io_in_stage(local_pes_21_8_io_in_stage),
    .io_out_q(local_pes_21_8_io_out_q),
    .io_out_sum(local_pes_21_8_io_out_sum),
    .io_out_sum_exp(local_pes_21_8_io_out_sum_exp),
    .io_out_kv(local_pes_21_8_io_out_kv),
    .io_out_stage(local_pes_21_8_io_out_stage)
  );
  PE_1 local_pes_21_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_9_clock),
    .reset(local_pes_21_9_reset),
    .io_in_q(local_pes_21_9_io_in_q),
    .io_in_sum(local_pes_21_9_io_in_sum),
    .io_in_sum_exp(local_pes_21_9_io_in_sum_exp),
    .io_in_kv(local_pes_21_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_9_io_in_inv_sum),
    .io_in_stage(local_pes_21_9_io_in_stage),
    .io_out_q(local_pes_21_9_io_out_q),
    .io_out_sum(local_pes_21_9_io_out_sum),
    .io_out_sum_exp(local_pes_21_9_io_out_sum_exp),
    .io_out_kv(local_pes_21_9_io_out_kv),
    .io_out_stage(local_pes_21_9_io_out_stage)
  );
  PE_1 local_pes_21_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_10_clock),
    .reset(local_pes_21_10_reset),
    .io_in_q(local_pes_21_10_io_in_q),
    .io_in_sum(local_pes_21_10_io_in_sum),
    .io_in_sum_exp(local_pes_21_10_io_in_sum_exp),
    .io_in_kv(local_pes_21_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_10_io_in_inv_sum),
    .io_in_stage(local_pes_21_10_io_in_stage),
    .io_out_q(local_pes_21_10_io_out_q),
    .io_out_sum(local_pes_21_10_io_out_sum),
    .io_out_sum_exp(local_pes_21_10_io_out_sum_exp),
    .io_out_kv(local_pes_21_10_io_out_kv),
    .io_out_stage(local_pes_21_10_io_out_stage)
  );
  PE_1 local_pes_21_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_11_clock),
    .reset(local_pes_21_11_reset),
    .io_in_q(local_pes_21_11_io_in_q),
    .io_in_sum(local_pes_21_11_io_in_sum),
    .io_in_sum_exp(local_pes_21_11_io_in_sum_exp),
    .io_in_kv(local_pes_21_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_11_io_in_inv_sum),
    .io_in_stage(local_pes_21_11_io_in_stage),
    .io_out_q(local_pes_21_11_io_out_q),
    .io_out_sum(local_pes_21_11_io_out_sum),
    .io_out_sum_exp(local_pes_21_11_io_out_sum_exp),
    .io_out_kv(local_pes_21_11_io_out_kv),
    .io_out_stage(local_pes_21_11_io_out_stage)
  );
  PE_1 local_pes_21_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_12_clock),
    .reset(local_pes_21_12_reset),
    .io_in_q(local_pes_21_12_io_in_q),
    .io_in_sum(local_pes_21_12_io_in_sum),
    .io_in_sum_exp(local_pes_21_12_io_in_sum_exp),
    .io_in_kv(local_pes_21_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_12_io_in_inv_sum),
    .io_in_stage(local_pes_21_12_io_in_stage),
    .io_out_q(local_pes_21_12_io_out_q),
    .io_out_sum(local_pes_21_12_io_out_sum),
    .io_out_sum_exp(local_pes_21_12_io_out_sum_exp),
    .io_out_kv(local_pes_21_12_io_out_kv),
    .io_out_stage(local_pes_21_12_io_out_stage)
  );
  PE_1 local_pes_21_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_13_clock),
    .reset(local_pes_21_13_reset),
    .io_in_q(local_pes_21_13_io_in_q),
    .io_in_sum(local_pes_21_13_io_in_sum),
    .io_in_sum_exp(local_pes_21_13_io_in_sum_exp),
    .io_in_kv(local_pes_21_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_13_io_in_inv_sum),
    .io_in_stage(local_pes_21_13_io_in_stage),
    .io_out_q(local_pes_21_13_io_out_q),
    .io_out_sum(local_pes_21_13_io_out_sum),
    .io_out_sum_exp(local_pes_21_13_io_out_sum_exp),
    .io_out_kv(local_pes_21_13_io_out_kv),
    .io_out_stage(local_pes_21_13_io_out_stage)
  );
  PE_1 local_pes_21_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_14_clock),
    .reset(local_pes_21_14_reset),
    .io_in_q(local_pes_21_14_io_in_q),
    .io_in_sum(local_pes_21_14_io_in_sum),
    .io_in_sum_exp(local_pes_21_14_io_in_sum_exp),
    .io_in_kv(local_pes_21_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_14_io_in_inv_sum),
    .io_in_stage(local_pes_21_14_io_in_stage),
    .io_out_q(local_pes_21_14_io_out_q),
    .io_out_sum(local_pes_21_14_io_out_sum),
    .io_out_sum_exp(local_pes_21_14_io_out_sum_exp),
    .io_out_kv(local_pes_21_14_io_out_kv),
    .io_out_stage(local_pes_21_14_io_out_stage)
  );
  PE_1 local_pes_21_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_15_clock),
    .reset(local_pes_21_15_reset),
    .io_in_q(local_pes_21_15_io_in_q),
    .io_in_sum(local_pes_21_15_io_in_sum),
    .io_in_sum_exp(local_pes_21_15_io_in_sum_exp),
    .io_in_kv(local_pes_21_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_15_io_in_inv_sum),
    .io_in_stage(local_pes_21_15_io_in_stage),
    .io_out_q(local_pes_21_15_io_out_q),
    .io_out_sum(local_pes_21_15_io_out_sum),
    .io_out_sum_exp(local_pes_21_15_io_out_sum_exp),
    .io_out_kv(local_pes_21_15_io_out_kv),
    .io_out_stage(local_pes_21_15_io_out_stage)
  );
  PE_1 local_pes_21_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_16_clock),
    .reset(local_pes_21_16_reset),
    .io_in_q(local_pes_21_16_io_in_q),
    .io_in_sum(local_pes_21_16_io_in_sum),
    .io_in_sum_exp(local_pes_21_16_io_in_sum_exp),
    .io_in_kv(local_pes_21_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_16_io_in_inv_sum),
    .io_in_stage(local_pes_21_16_io_in_stage),
    .io_out_q(local_pes_21_16_io_out_q),
    .io_out_sum(local_pes_21_16_io_out_sum),
    .io_out_sum_exp(local_pes_21_16_io_out_sum_exp),
    .io_out_kv(local_pes_21_16_io_out_kv),
    .io_out_stage(local_pes_21_16_io_out_stage)
  );
  PE_1 local_pes_21_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_17_clock),
    .reset(local_pes_21_17_reset),
    .io_in_q(local_pes_21_17_io_in_q),
    .io_in_sum(local_pes_21_17_io_in_sum),
    .io_in_sum_exp(local_pes_21_17_io_in_sum_exp),
    .io_in_kv(local_pes_21_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_17_io_in_inv_sum),
    .io_in_stage(local_pes_21_17_io_in_stage),
    .io_out_q(local_pes_21_17_io_out_q),
    .io_out_sum(local_pes_21_17_io_out_sum),
    .io_out_sum_exp(local_pes_21_17_io_out_sum_exp),
    .io_out_kv(local_pes_21_17_io_out_kv),
    .io_out_stage(local_pes_21_17_io_out_stage)
  );
  PE_1 local_pes_21_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_18_clock),
    .reset(local_pes_21_18_reset),
    .io_in_q(local_pes_21_18_io_in_q),
    .io_in_sum(local_pes_21_18_io_in_sum),
    .io_in_sum_exp(local_pes_21_18_io_in_sum_exp),
    .io_in_kv(local_pes_21_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_18_io_in_inv_sum),
    .io_in_stage(local_pes_21_18_io_in_stage),
    .io_out_q(local_pes_21_18_io_out_q),
    .io_out_sum(local_pes_21_18_io_out_sum),
    .io_out_sum_exp(local_pes_21_18_io_out_sum_exp),
    .io_out_kv(local_pes_21_18_io_out_kv),
    .io_out_stage(local_pes_21_18_io_out_stage)
  );
  PE_1 local_pes_21_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_19_clock),
    .reset(local_pes_21_19_reset),
    .io_in_q(local_pes_21_19_io_in_q),
    .io_in_sum(local_pes_21_19_io_in_sum),
    .io_in_sum_exp(local_pes_21_19_io_in_sum_exp),
    .io_in_kv(local_pes_21_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_19_io_in_inv_sum),
    .io_in_stage(local_pes_21_19_io_in_stage),
    .io_out_q(local_pes_21_19_io_out_q),
    .io_out_sum(local_pes_21_19_io_out_sum),
    .io_out_sum_exp(local_pes_21_19_io_out_sum_exp),
    .io_out_kv(local_pes_21_19_io_out_kv),
    .io_out_stage(local_pes_21_19_io_out_stage)
  );
  PE_1 local_pes_21_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_20_clock),
    .reset(local_pes_21_20_reset),
    .io_in_q(local_pes_21_20_io_in_q),
    .io_in_sum(local_pes_21_20_io_in_sum),
    .io_in_sum_exp(local_pes_21_20_io_in_sum_exp),
    .io_in_kv(local_pes_21_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_20_io_in_inv_sum),
    .io_in_stage(local_pes_21_20_io_in_stage),
    .io_out_q(local_pes_21_20_io_out_q),
    .io_out_sum(local_pes_21_20_io_out_sum),
    .io_out_sum_exp(local_pes_21_20_io_out_sum_exp),
    .io_out_kv(local_pes_21_20_io_out_kv),
    .io_out_stage(local_pes_21_20_io_out_stage)
  );
  PE_1 local_pes_21_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_21_clock),
    .reset(local_pes_21_21_reset),
    .io_in_q(local_pes_21_21_io_in_q),
    .io_in_sum(local_pes_21_21_io_in_sum),
    .io_in_sum_exp(local_pes_21_21_io_in_sum_exp),
    .io_in_kv(local_pes_21_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_21_io_in_inv_sum),
    .io_in_stage(local_pes_21_21_io_in_stage),
    .io_out_q(local_pes_21_21_io_out_q),
    .io_out_sum(local_pes_21_21_io_out_sum),
    .io_out_sum_exp(local_pes_21_21_io_out_sum_exp),
    .io_out_kv(local_pes_21_21_io_out_kv),
    .io_out_stage(local_pes_21_21_io_out_stage)
  );
  PE_1 local_pes_21_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_22_clock),
    .reset(local_pes_21_22_reset),
    .io_in_q(local_pes_21_22_io_in_q),
    .io_in_sum(local_pes_21_22_io_in_sum),
    .io_in_sum_exp(local_pes_21_22_io_in_sum_exp),
    .io_in_kv(local_pes_21_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_22_io_in_inv_sum),
    .io_in_stage(local_pes_21_22_io_in_stage),
    .io_out_q(local_pes_21_22_io_out_q),
    .io_out_sum(local_pes_21_22_io_out_sum),
    .io_out_sum_exp(local_pes_21_22_io_out_sum_exp),
    .io_out_kv(local_pes_21_22_io_out_kv),
    .io_out_stage(local_pes_21_22_io_out_stage)
  );
  PE_1 local_pes_21_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_23_clock),
    .reset(local_pes_21_23_reset),
    .io_in_q(local_pes_21_23_io_in_q),
    .io_in_sum(local_pes_21_23_io_in_sum),
    .io_in_sum_exp(local_pes_21_23_io_in_sum_exp),
    .io_in_kv(local_pes_21_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_23_io_in_inv_sum),
    .io_in_stage(local_pes_21_23_io_in_stage),
    .io_out_q(local_pes_21_23_io_out_q),
    .io_out_sum(local_pes_21_23_io_out_sum),
    .io_out_sum_exp(local_pes_21_23_io_out_sum_exp),
    .io_out_kv(local_pes_21_23_io_out_kv),
    .io_out_stage(local_pes_21_23_io_out_stage)
  );
  PE_1 local_pes_21_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_24_clock),
    .reset(local_pes_21_24_reset),
    .io_in_q(local_pes_21_24_io_in_q),
    .io_in_sum(local_pes_21_24_io_in_sum),
    .io_in_sum_exp(local_pes_21_24_io_in_sum_exp),
    .io_in_kv(local_pes_21_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_24_io_in_inv_sum),
    .io_in_stage(local_pes_21_24_io_in_stage),
    .io_out_q(local_pes_21_24_io_out_q),
    .io_out_sum(local_pes_21_24_io_out_sum),
    .io_out_sum_exp(local_pes_21_24_io_out_sum_exp),
    .io_out_kv(local_pes_21_24_io_out_kv),
    .io_out_stage(local_pes_21_24_io_out_stage)
  );
  PE_1 local_pes_21_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_25_clock),
    .reset(local_pes_21_25_reset),
    .io_in_q(local_pes_21_25_io_in_q),
    .io_in_sum(local_pes_21_25_io_in_sum),
    .io_in_sum_exp(local_pes_21_25_io_in_sum_exp),
    .io_in_kv(local_pes_21_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_25_io_in_inv_sum),
    .io_in_stage(local_pes_21_25_io_in_stage),
    .io_out_q(local_pes_21_25_io_out_q),
    .io_out_sum(local_pes_21_25_io_out_sum),
    .io_out_sum_exp(local_pes_21_25_io_out_sum_exp),
    .io_out_kv(local_pes_21_25_io_out_kv),
    .io_out_stage(local_pes_21_25_io_out_stage)
  );
  PE_1 local_pes_21_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_26_clock),
    .reset(local_pes_21_26_reset),
    .io_in_q(local_pes_21_26_io_in_q),
    .io_in_sum(local_pes_21_26_io_in_sum),
    .io_in_sum_exp(local_pes_21_26_io_in_sum_exp),
    .io_in_kv(local_pes_21_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_26_io_in_inv_sum),
    .io_in_stage(local_pes_21_26_io_in_stage),
    .io_out_q(local_pes_21_26_io_out_q),
    .io_out_sum(local_pes_21_26_io_out_sum),
    .io_out_sum_exp(local_pes_21_26_io_out_sum_exp),
    .io_out_kv(local_pes_21_26_io_out_kv),
    .io_out_stage(local_pes_21_26_io_out_stage)
  );
  PE_1 local_pes_21_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_27_clock),
    .reset(local_pes_21_27_reset),
    .io_in_q(local_pes_21_27_io_in_q),
    .io_in_sum(local_pes_21_27_io_in_sum),
    .io_in_sum_exp(local_pes_21_27_io_in_sum_exp),
    .io_in_kv(local_pes_21_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_27_io_in_inv_sum),
    .io_in_stage(local_pes_21_27_io_in_stage),
    .io_out_q(local_pes_21_27_io_out_q),
    .io_out_sum(local_pes_21_27_io_out_sum),
    .io_out_sum_exp(local_pes_21_27_io_out_sum_exp),
    .io_out_kv(local_pes_21_27_io_out_kv),
    .io_out_stage(local_pes_21_27_io_out_stage)
  );
  PE_1 local_pes_21_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_28_clock),
    .reset(local_pes_21_28_reset),
    .io_in_q(local_pes_21_28_io_in_q),
    .io_in_sum(local_pes_21_28_io_in_sum),
    .io_in_sum_exp(local_pes_21_28_io_in_sum_exp),
    .io_in_kv(local_pes_21_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_28_io_in_inv_sum),
    .io_in_stage(local_pes_21_28_io_in_stage),
    .io_out_q(local_pes_21_28_io_out_q),
    .io_out_sum(local_pes_21_28_io_out_sum),
    .io_out_sum_exp(local_pes_21_28_io_out_sum_exp),
    .io_out_kv(local_pes_21_28_io_out_kv),
    .io_out_stage(local_pes_21_28_io_out_stage)
  );
  PE_1 local_pes_21_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_29_clock),
    .reset(local_pes_21_29_reset),
    .io_in_q(local_pes_21_29_io_in_q),
    .io_in_sum(local_pes_21_29_io_in_sum),
    .io_in_sum_exp(local_pes_21_29_io_in_sum_exp),
    .io_in_kv(local_pes_21_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_29_io_in_inv_sum),
    .io_in_stage(local_pes_21_29_io_in_stage),
    .io_out_q(local_pes_21_29_io_out_q),
    .io_out_sum(local_pes_21_29_io_out_sum),
    .io_out_sum_exp(local_pes_21_29_io_out_sum_exp),
    .io_out_kv(local_pes_21_29_io_out_kv),
    .io_out_stage(local_pes_21_29_io_out_stage)
  );
  PE_1 local_pes_21_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_30_clock),
    .reset(local_pes_21_30_reset),
    .io_in_q(local_pes_21_30_io_in_q),
    .io_in_sum(local_pes_21_30_io_in_sum),
    .io_in_sum_exp(local_pes_21_30_io_in_sum_exp),
    .io_in_kv(local_pes_21_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_30_io_in_inv_sum),
    .io_in_stage(local_pes_21_30_io_in_stage),
    .io_out_q(local_pes_21_30_io_out_q),
    .io_out_sum(local_pes_21_30_io_out_sum),
    .io_out_sum_exp(local_pes_21_30_io_out_sum_exp),
    .io_out_kv(local_pes_21_30_io_out_kv),
    .io_out_stage(local_pes_21_30_io_out_stage)
  );
  PE_1 local_pes_21_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_21_31_clock),
    .reset(local_pes_21_31_reset),
    .io_in_q(local_pes_21_31_io_in_q),
    .io_in_sum(local_pes_21_31_io_in_sum),
    .io_in_sum_exp(local_pes_21_31_io_in_sum_exp),
    .io_in_kv(local_pes_21_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_21_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_21_31_io_in_inv_sum),
    .io_in_stage(local_pes_21_31_io_in_stage),
    .io_out_q(local_pes_21_31_io_out_q),
    .io_out_sum(local_pes_21_31_io_out_sum),
    .io_out_sum_exp(local_pes_21_31_io_out_sum_exp),
    .io_out_kv(local_pes_21_31_io_out_kv),
    .io_out_stage(local_pes_21_31_io_out_stage)
  );
  PE local_pes_22_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_0_clock),
    .reset(local_pes_22_0_reset),
    .io_in_q(local_pes_22_0_io_in_q),
    .io_in_kv(local_pes_22_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_0_io_in_inv_sum),
    .io_in_stage(local_pes_22_0_io_in_stage),
    .io_out_q(local_pes_22_0_io_out_q),
    .io_out_sum(local_pes_22_0_io_out_sum),
    .io_out_kv(local_pes_22_0_io_out_kv),
    .io_out_stage(local_pes_22_0_io_out_stage)
  );
  PE_1 local_pes_22_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_1_clock),
    .reset(local_pes_22_1_reset),
    .io_in_q(local_pes_22_1_io_in_q),
    .io_in_sum(local_pes_22_1_io_in_sum),
    .io_in_sum_exp(local_pes_22_1_io_in_sum_exp),
    .io_in_kv(local_pes_22_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_1_io_in_inv_sum),
    .io_in_stage(local_pes_22_1_io_in_stage),
    .io_out_q(local_pes_22_1_io_out_q),
    .io_out_sum(local_pes_22_1_io_out_sum),
    .io_out_sum_exp(local_pes_22_1_io_out_sum_exp),
    .io_out_kv(local_pes_22_1_io_out_kv),
    .io_out_stage(local_pes_22_1_io_out_stage)
  );
  PE_1 local_pes_22_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_2_clock),
    .reset(local_pes_22_2_reset),
    .io_in_q(local_pes_22_2_io_in_q),
    .io_in_sum(local_pes_22_2_io_in_sum),
    .io_in_sum_exp(local_pes_22_2_io_in_sum_exp),
    .io_in_kv(local_pes_22_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_2_io_in_inv_sum),
    .io_in_stage(local_pes_22_2_io_in_stage),
    .io_out_q(local_pes_22_2_io_out_q),
    .io_out_sum(local_pes_22_2_io_out_sum),
    .io_out_sum_exp(local_pes_22_2_io_out_sum_exp),
    .io_out_kv(local_pes_22_2_io_out_kv),
    .io_out_stage(local_pes_22_2_io_out_stage)
  );
  PE_1 local_pes_22_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_3_clock),
    .reset(local_pes_22_3_reset),
    .io_in_q(local_pes_22_3_io_in_q),
    .io_in_sum(local_pes_22_3_io_in_sum),
    .io_in_sum_exp(local_pes_22_3_io_in_sum_exp),
    .io_in_kv(local_pes_22_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_3_io_in_inv_sum),
    .io_in_stage(local_pes_22_3_io_in_stage),
    .io_out_q(local_pes_22_3_io_out_q),
    .io_out_sum(local_pes_22_3_io_out_sum),
    .io_out_sum_exp(local_pes_22_3_io_out_sum_exp),
    .io_out_kv(local_pes_22_3_io_out_kv),
    .io_out_stage(local_pes_22_3_io_out_stage)
  );
  PE_1 local_pes_22_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_4_clock),
    .reset(local_pes_22_4_reset),
    .io_in_q(local_pes_22_4_io_in_q),
    .io_in_sum(local_pes_22_4_io_in_sum),
    .io_in_sum_exp(local_pes_22_4_io_in_sum_exp),
    .io_in_kv(local_pes_22_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_4_io_in_inv_sum),
    .io_in_stage(local_pes_22_4_io_in_stage),
    .io_out_q(local_pes_22_4_io_out_q),
    .io_out_sum(local_pes_22_4_io_out_sum),
    .io_out_sum_exp(local_pes_22_4_io_out_sum_exp),
    .io_out_kv(local_pes_22_4_io_out_kv),
    .io_out_stage(local_pes_22_4_io_out_stage)
  );
  PE_1 local_pes_22_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_5_clock),
    .reset(local_pes_22_5_reset),
    .io_in_q(local_pes_22_5_io_in_q),
    .io_in_sum(local_pes_22_5_io_in_sum),
    .io_in_sum_exp(local_pes_22_5_io_in_sum_exp),
    .io_in_kv(local_pes_22_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_5_io_in_inv_sum),
    .io_in_stage(local_pes_22_5_io_in_stage),
    .io_out_q(local_pes_22_5_io_out_q),
    .io_out_sum(local_pes_22_5_io_out_sum),
    .io_out_sum_exp(local_pes_22_5_io_out_sum_exp),
    .io_out_kv(local_pes_22_5_io_out_kv),
    .io_out_stage(local_pes_22_5_io_out_stage)
  );
  PE_1 local_pes_22_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_6_clock),
    .reset(local_pes_22_6_reset),
    .io_in_q(local_pes_22_6_io_in_q),
    .io_in_sum(local_pes_22_6_io_in_sum),
    .io_in_sum_exp(local_pes_22_6_io_in_sum_exp),
    .io_in_kv(local_pes_22_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_6_io_in_inv_sum),
    .io_in_stage(local_pes_22_6_io_in_stage),
    .io_out_q(local_pes_22_6_io_out_q),
    .io_out_sum(local_pes_22_6_io_out_sum),
    .io_out_sum_exp(local_pes_22_6_io_out_sum_exp),
    .io_out_kv(local_pes_22_6_io_out_kv),
    .io_out_stage(local_pes_22_6_io_out_stage)
  );
  PE_1 local_pes_22_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_7_clock),
    .reset(local_pes_22_7_reset),
    .io_in_q(local_pes_22_7_io_in_q),
    .io_in_sum(local_pes_22_7_io_in_sum),
    .io_in_sum_exp(local_pes_22_7_io_in_sum_exp),
    .io_in_kv(local_pes_22_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_7_io_in_inv_sum),
    .io_in_stage(local_pes_22_7_io_in_stage),
    .io_out_q(local_pes_22_7_io_out_q),
    .io_out_sum(local_pes_22_7_io_out_sum),
    .io_out_sum_exp(local_pes_22_7_io_out_sum_exp),
    .io_out_kv(local_pes_22_7_io_out_kv),
    .io_out_stage(local_pes_22_7_io_out_stage)
  );
  PE_1 local_pes_22_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_8_clock),
    .reset(local_pes_22_8_reset),
    .io_in_q(local_pes_22_8_io_in_q),
    .io_in_sum(local_pes_22_8_io_in_sum),
    .io_in_sum_exp(local_pes_22_8_io_in_sum_exp),
    .io_in_kv(local_pes_22_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_8_io_in_inv_sum),
    .io_in_stage(local_pes_22_8_io_in_stage),
    .io_out_q(local_pes_22_8_io_out_q),
    .io_out_sum(local_pes_22_8_io_out_sum),
    .io_out_sum_exp(local_pes_22_8_io_out_sum_exp),
    .io_out_kv(local_pes_22_8_io_out_kv),
    .io_out_stage(local_pes_22_8_io_out_stage)
  );
  PE_1 local_pes_22_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_9_clock),
    .reset(local_pes_22_9_reset),
    .io_in_q(local_pes_22_9_io_in_q),
    .io_in_sum(local_pes_22_9_io_in_sum),
    .io_in_sum_exp(local_pes_22_9_io_in_sum_exp),
    .io_in_kv(local_pes_22_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_9_io_in_inv_sum),
    .io_in_stage(local_pes_22_9_io_in_stage),
    .io_out_q(local_pes_22_9_io_out_q),
    .io_out_sum(local_pes_22_9_io_out_sum),
    .io_out_sum_exp(local_pes_22_9_io_out_sum_exp),
    .io_out_kv(local_pes_22_9_io_out_kv),
    .io_out_stage(local_pes_22_9_io_out_stage)
  );
  PE_1 local_pes_22_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_10_clock),
    .reset(local_pes_22_10_reset),
    .io_in_q(local_pes_22_10_io_in_q),
    .io_in_sum(local_pes_22_10_io_in_sum),
    .io_in_sum_exp(local_pes_22_10_io_in_sum_exp),
    .io_in_kv(local_pes_22_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_10_io_in_inv_sum),
    .io_in_stage(local_pes_22_10_io_in_stage),
    .io_out_q(local_pes_22_10_io_out_q),
    .io_out_sum(local_pes_22_10_io_out_sum),
    .io_out_sum_exp(local_pes_22_10_io_out_sum_exp),
    .io_out_kv(local_pes_22_10_io_out_kv),
    .io_out_stage(local_pes_22_10_io_out_stage)
  );
  PE_1 local_pes_22_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_11_clock),
    .reset(local_pes_22_11_reset),
    .io_in_q(local_pes_22_11_io_in_q),
    .io_in_sum(local_pes_22_11_io_in_sum),
    .io_in_sum_exp(local_pes_22_11_io_in_sum_exp),
    .io_in_kv(local_pes_22_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_11_io_in_inv_sum),
    .io_in_stage(local_pes_22_11_io_in_stage),
    .io_out_q(local_pes_22_11_io_out_q),
    .io_out_sum(local_pes_22_11_io_out_sum),
    .io_out_sum_exp(local_pes_22_11_io_out_sum_exp),
    .io_out_kv(local_pes_22_11_io_out_kv),
    .io_out_stage(local_pes_22_11_io_out_stage)
  );
  PE_1 local_pes_22_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_12_clock),
    .reset(local_pes_22_12_reset),
    .io_in_q(local_pes_22_12_io_in_q),
    .io_in_sum(local_pes_22_12_io_in_sum),
    .io_in_sum_exp(local_pes_22_12_io_in_sum_exp),
    .io_in_kv(local_pes_22_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_12_io_in_inv_sum),
    .io_in_stage(local_pes_22_12_io_in_stage),
    .io_out_q(local_pes_22_12_io_out_q),
    .io_out_sum(local_pes_22_12_io_out_sum),
    .io_out_sum_exp(local_pes_22_12_io_out_sum_exp),
    .io_out_kv(local_pes_22_12_io_out_kv),
    .io_out_stage(local_pes_22_12_io_out_stage)
  );
  PE_1 local_pes_22_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_13_clock),
    .reset(local_pes_22_13_reset),
    .io_in_q(local_pes_22_13_io_in_q),
    .io_in_sum(local_pes_22_13_io_in_sum),
    .io_in_sum_exp(local_pes_22_13_io_in_sum_exp),
    .io_in_kv(local_pes_22_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_13_io_in_inv_sum),
    .io_in_stage(local_pes_22_13_io_in_stage),
    .io_out_q(local_pes_22_13_io_out_q),
    .io_out_sum(local_pes_22_13_io_out_sum),
    .io_out_sum_exp(local_pes_22_13_io_out_sum_exp),
    .io_out_kv(local_pes_22_13_io_out_kv),
    .io_out_stage(local_pes_22_13_io_out_stage)
  );
  PE_1 local_pes_22_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_14_clock),
    .reset(local_pes_22_14_reset),
    .io_in_q(local_pes_22_14_io_in_q),
    .io_in_sum(local_pes_22_14_io_in_sum),
    .io_in_sum_exp(local_pes_22_14_io_in_sum_exp),
    .io_in_kv(local_pes_22_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_14_io_in_inv_sum),
    .io_in_stage(local_pes_22_14_io_in_stage),
    .io_out_q(local_pes_22_14_io_out_q),
    .io_out_sum(local_pes_22_14_io_out_sum),
    .io_out_sum_exp(local_pes_22_14_io_out_sum_exp),
    .io_out_kv(local_pes_22_14_io_out_kv),
    .io_out_stage(local_pes_22_14_io_out_stage)
  );
  PE_1 local_pes_22_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_15_clock),
    .reset(local_pes_22_15_reset),
    .io_in_q(local_pes_22_15_io_in_q),
    .io_in_sum(local_pes_22_15_io_in_sum),
    .io_in_sum_exp(local_pes_22_15_io_in_sum_exp),
    .io_in_kv(local_pes_22_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_15_io_in_inv_sum),
    .io_in_stage(local_pes_22_15_io_in_stage),
    .io_out_q(local_pes_22_15_io_out_q),
    .io_out_sum(local_pes_22_15_io_out_sum),
    .io_out_sum_exp(local_pes_22_15_io_out_sum_exp),
    .io_out_kv(local_pes_22_15_io_out_kv),
    .io_out_stage(local_pes_22_15_io_out_stage)
  );
  PE_1 local_pes_22_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_16_clock),
    .reset(local_pes_22_16_reset),
    .io_in_q(local_pes_22_16_io_in_q),
    .io_in_sum(local_pes_22_16_io_in_sum),
    .io_in_sum_exp(local_pes_22_16_io_in_sum_exp),
    .io_in_kv(local_pes_22_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_16_io_in_inv_sum),
    .io_in_stage(local_pes_22_16_io_in_stage),
    .io_out_q(local_pes_22_16_io_out_q),
    .io_out_sum(local_pes_22_16_io_out_sum),
    .io_out_sum_exp(local_pes_22_16_io_out_sum_exp),
    .io_out_kv(local_pes_22_16_io_out_kv),
    .io_out_stage(local_pes_22_16_io_out_stage)
  );
  PE_1 local_pes_22_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_17_clock),
    .reset(local_pes_22_17_reset),
    .io_in_q(local_pes_22_17_io_in_q),
    .io_in_sum(local_pes_22_17_io_in_sum),
    .io_in_sum_exp(local_pes_22_17_io_in_sum_exp),
    .io_in_kv(local_pes_22_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_17_io_in_inv_sum),
    .io_in_stage(local_pes_22_17_io_in_stage),
    .io_out_q(local_pes_22_17_io_out_q),
    .io_out_sum(local_pes_22_17_io_out_sum),
    .io_out_sum_exp(local_pes_22_17_io_out_sum_exp),
    .io_out_kv(local_pes_22_17_io_out_kv),
    .io_out_stage(local_pes_22_17_io_out_stage)
  );
  PE_1 local_pes_22_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_18_clock),
    .reset(local_pes_22_18_reset),
    .io_in_q(local_pes_22_18_io_in_q),
    .io_in_sum(local_pes_22_18_io_in_sum),
    .io_in_sum_exp(local_pes_22_18_io_in_sum_exp),
    .io_in_kv(local_pes_22_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_18_io_in_inv_sum),
    .io_in_stage(local_pes_22_18_io_in_stage),
    .io_out_q(local_pes_22_18_io_out_q),
    .io_out_sum(local_pes_22_18_io_out_sum),
    .io_out_sum_exp(local_pes_22_18_io_out_sum_exp),
    .io_out_kv(local_pes_22_18_io_out_kv),
    .io_out_stage(local_pes_22_18_io_out_stage)
  );
  PE_1 local_pes_22_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_19_clock),
    .reset(local_pes_22_19_reset),
    .io_in_q(local_pes_22_19_io_in_q),
    .io_in_sum(local_pes_22_19_io_in_sum),
    .io_in_sum_exp(local_pes_22_19_io_in_sum_exp),
    .io_in_kv(local_pes_22_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_19_io_in_inv_sum),
    .io_in_stage(local_pes_22_19_io_in_stage),
    .io_out_q(local_pes_22_19_io_out_q),
    .io_out_sum(local_pes_22_19_io_out_sum),
    .io_out_sum_exp(local_pes_22_19_io_out_sum_exp),
    .io_out_kv(local_pes_22_19_io_out_kv),
    .io_out_stage(local_pes_22_19_io_out_stage)
  );
  PE_1 local_pes_22_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_20_clock),
    .reset(local_pes_22_20_reset),
    .io_in_q(local_pes_22_20_io_in_q),
    .io_in_sum(local_pes_22_20_io_in_sum),
    .io_in_sum_exp(local_pes_22_20_io_in_sum_exp),
    .io_in_kv(local_pes_22_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_20_io_in_inv_sum),
    .io_in_stage(local_pes_22_20_io_in_stage),
    .io_out_q(local_pes_22_20_io_out_q),
    .io_out_sum(local_pes_22_20_io_out_sum),
    .io_out_sum_exp(local_pes_22_20_io_out_sum_exp),
    .io_out_kv(local_pes_22_20_io_out_kv),
    .io_out_stage(local_pes_22_20_io_out_stage)
  );
  PE_1 local_pes_22_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_21_clock),
    .reset(local_pes_22_21_reset),
    .io_in_q(local_pes_22_21_io_in_q),
    .io_in_sum(local_pes_22_21_io_in_sum),
    .io_in_sum_exp(local_pes_22_21_io_in_sum_exp),
    .io_in_kv(local_pes_22_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_21_io_in_inv_sum),
    .io_in_stage(local_pes_22_21_io_in_stage),
    .io_out_q(local_pes_22_21_io_out_q),
    .io_out_sum(local_pes_22_21_io_out_sum),
    .io_out_sum_exp(local_pes_22_21_io_out_sum_exp),
    .io_out_kv(local_pes_22_21_io_out_kv),
    .io_out_stage(local_pes_22_21_io_out_stage)
  );
  PE_1 local_pes_22_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_22_clock),
    .reset(local_pes_22_22_reset),
    .io_in_q(local_pes_22_22_io_in_q),
    .io_in_sum(local_pes_22_22_io_in_sum),
    .io_in_sum_exp(local_pes_22_22_io_in_sum_exp),
    .io_in_kv(local_pes_22_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_22_io_in_inv_sum),
    .io_in_stage(local_pes_22_22_io_in_stage),
    .io_out_q(local_pes_22_22_io_out_q),
    .io_out_sum(local_pes_22_22_io_out_sum),
    .io_out_sum_exp(local_pes_22_22_io_out_sum_exp),
    .io_out_kv(local_pes_22_22_io_out_kv),
    .io_out_stage(local_pes_22_22_io_out_stage)
  );
  PE_1 local_pes_22_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_23_clock),
    .reset(local_pes_22_23_reset),
    .io_in_q(local_pes_22_23_io_in_q),
    .io_in_sum(local_pes_22_23_io_in_sum),
    .io_in_sum_exp(local_pes_22_23_io_in_sum_exp),
    .io_in_kv(local_pes_22_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_23_io_in_inv_sum),
    .io_in_stage(local_pes_22_23_io_in_stage),
    .io_out_q(local_pes_22_23_io_out_q),
    .io_out_sum(local_pes_22_23_io_out_sum),
    .io_out_sum_exp(local_pes_22_23_io_out_sum_exp),
    .io_out_kv(local_pes_22_23_io_out_kv),
    .io_out_stage(local_pes_22_23_io_out_stage)
  );
  PE_1 local_pes_22_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_24_clock),
    .reset(local_pes_22_24_reset),
    .io_in_q(local_pes_22_24_io_in_q),
    .io_in_sum(local_pes_22_24_io_in_sum),
    .io_in_sum_exp(local_pes_22_24_io_in_sum_exp),
    .io_in_kv(local_pes_22_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_24_io_in_inv_sum),
    .io_in_stage(local_pes_22_24_io_in_stage),
    .io_out_q(local_pes_22_24_io_out_q),
    .io_out_sum(local_pes_22_24_io_out_sum),
    .io_out_sum_exp(local_pes_22_24_io_out_sum_exp),
    .io_out_kv(local_pes_22_24_io_out_kv),
    .io_out_stage(local_pes_22_24_io_out_stage)
  );
  PE_1 local_pes_22_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_25_clock),
    .reset(local_pes_22_25_reset),
    .io_in_q(local_pes_22_25_io_in_q),
    .io_in_sum(local_pes_22_25_io_in_sum),
    .io_in_sum_exp(local_pes_22_25_io_in_sum_exp),
    .io_in_kv(local_pes_22_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_25_io_in_inv_sum),
    .io_in_stage(local_pes_22_25_io_in_stage),
    .io_out_q(local_pes_22_25_io_out_q),
    .io_out_sum(local_pes_22_25_io_out_sum),
    .io_out_sum_exp(local_pes_22_25_io_out_sum_exp),
    .io_out_kv(local_pes_22_25_io_out_kv),
    .io_out_stage(local_pes_22_25_io_out_stage)
  );
  PE_1 local_pes_22_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_26_clock),
    .reset(local_pes_22_26_reset),
    .io_in_q(local_pes_22_26_io_in_q),
    .io_in_sum(local_pes_22_26_io_in_sum),
    .io_in_sum_exp(local_pes_22_26_io_in_sum_exp),
    .io_in_kv(local_pes_22_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_26_io_in_inv_sum),
    .io_in_stage(local_pes_22_26_io_in_stage),
    .io_out_q(local_pes_22_26_io_out_q),
    .io_out_sum(local_pes_22_26_io_out_sum),
    .io_out_sum_exp(local_pes_22_26_io_out_sum_exp),
    .io_out_kv(local_pes_22_26_io_out_kv),
    .io_out_stage(local_pes_22_26_io_out_stage)
  );
  PE_1 local_pes_22_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_27_clock),
    .reset(local_pes_22_27_reset),
    .io_in_q(local_pes_22_27_io_in_q),
    .io_in_sum(local_pes_22_27_io_in_sum),
    .io_in_sum_exp(local_pes_22_27_io_in_sum_exp),
    .io_in_kv(local_pes_22_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_27_io_in_inv_sum),
    .io_in_stage(local_pes_22_27_io_in_stage),
    .io_out_q(local_pes_22_27_io_out_q),
    .io_out_sum(local_pes_22_27_io_out_sum),
    .io_out_sum_exp(local_pes_22_27_io_out_sum_exp),
    .io_out_kv(local_pes_22_27_io_out_kv),
    .io_out_stage(local_pes_22_27_io_out_stage)
  );
  PE_1 local_pes_22_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_28_clock),
    .reset(local_pes_22_28_reset),
    .io_in_q(local_pes_22_28_io_in_q),
    .io_in_sum(local_pes_22_28_io_in_sum),
    .io_in_sum_exp(local_pes_22_28_io_in_sum_exp),
    .io_in_kv(local_pes_22_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_28_io_in_inv_sum),
    .io_in_stage(local_pes_22_28_io_in_stage),
    .io_out_q(local_pes_22_28_io_out_q),
    .io_out_sum(local_pes_22_28_io_out_sum),
    .io_out_sum_exp(local_pes_22_28_io_out_sum_exp),
    .io_out_kv(local_pes_22_28_io_out_kv),
    .io_out_stage(local_pes_22_28_io_out_stage)
  );
  PE_1 local_pes_22_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_29_clock),
    .reset(local_pes_22_29_reset),
    .io_in_q(local_pes_22_29_io_in_q),
    .io_in_sum(local_pes_22_29_io_in_sum),
    .io_in_sum_exp(local_pes_22_29_io_in_sum_exp),
    .io_in_kv(local_pes_22_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_29_io_in_inv_sum),
    .io_in_stage(local_pes_22_29_io_in_stage),
    .io_out_q(local_pes_22_29_io_out_q),
    .io_out_sum(local_pes_22_29_io_out_sum),
    .io_out_sum_exp(local_pes_22_29_io_out_sum_exp),
    .io_out_kv(local_pes_22_29_io_out_kv),
    .io_out_stage(local_pes_22_29_io_out_stage)
  );
  PE_1 local_pes_22_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_30_clock),
    .reset(local_pes_22_30_reset),
    .io_in_q(local_pes_22_30_io_in_q),
    .io_in_sum(local_pes_22_30_io_in_sum),
    .io_in_sum_exp(local_pes_22_30_io_in_sum_exp),
    .io_in_kv(local_pes_22_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_30_io_in_inv_sum),
    .io_in_stage(local_pes_22_30_io_in_stage),
    .io_out_q(local_pes_22_30_io_out_q),
    .io_out_sum(local_pes_22_30_io_out_sum),
    .io_out_sum_exp(local_pes_22_30_io_out_sum_exp),
    .io_out_kv(local_pes_22_30_io_out_kv),
    .io_out_stage(local_pes_22_30_io_out_stage)
  );
  PE_1 local_pes_22_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_22_31_clock),
    .reset(local_pes_22_31_reset),
    .io_in_q(local_pes_22_31_io_in_q),
    .io_in_sum(local_pes_22_31_io_in_sum),
    .io_in_sum_exp(local_pes_22_31_io_in_sum_exp),
    .io_in_kv(local_pes_22_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_22_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_22_31_io_in_inv_sum),
    .io_in_stage(local_pes_22_31_io_in_stage),
    .io_out_q(local_pes_22_31_io_out_q),
    .io_out_sum(local_pes_22_31_io_out_sum),
    .io_out_sum_exp(local_pes_22_31_io_out_sum_exp),
    .io_out_kv(local_pes_22_31_io_out_kv),
    .io_out_stage(local_pes_22_31_io_out_stage)
  );
  PE local_pes_23_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_0_clock),
    .reset(local_pes_23_0_reset),
    .io_in_q(local_pes_23_0_io_in_q),
    .io_in_kv(local_pes_23_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_0_io_in_inv_sum),
    .io_in_stage(local_pes_23_0_io_in_stage),
    .io_out_q(local_pes_23_0_io_out_q),
    .io_out_sum(local_pes_23_0_io_out_sum),
    .io_out_kv(local_pes_23_0_io_out_kv),
    .io_out_stage(local_pes_23_0_io_out_stage)
  );
  PE_1 local_pes_23_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_1_clock),
    .reset(local_pes_23_1_reset),
    .io_in_q(local_pes_23_1_io_in_q),
    .io_in_sum(local_pes_23_1_io_in_sum),
    .io_in_sum_exp(local_pes_23_1_io_in_sum_exp),
    .io_in_kv(local_pes_23_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_1_io_in_inv_sum),
    .io_in_stage(local_pes_23_1_io_in_stage),
    .io_out_q(local_pes_23_1_io_out_q),
    .io_out_sum(local_pes_23_1_io_out_sum),
    .io_out_sum_exp(local_pes_23_1_io_out_sum_exp),
    .io_out_kv(local_pes_23_1_io_out_kv),
    .io_out_stage(local_pes_23_1_io_out_stage)
  );
  PE_1 local_pes_23_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_2_clock),
    .reset(local_pes_23_2_reset),
    .io_in_q(local_pes_23_2_io_in_q),
    .io_in_sum(local_pes_23_2_io_in_sum),
    .io_in_sum_exp(local_pes_23_2_io_in_sum_exp),
    .io_in_kv(local_pes_23_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_2_io_in_inv_sum),
    .io_in_stage(local_pes_23_2_io_in_stage),
    .io_out_q(local_pes_23_2_io_out_q),
    .io_out_sum(local_pes_23_2_io_out_sum),
    .io_out_sum_exp(local_pes_23_2_io_out_sum_exp),
    .io_out_kv(local_pes_23_2_io_out_kv),
    .io_out_stage(local_pes_23_2_io_out_stage)
  );
  PE_1 local_pes_23_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_3_clock),
    .reset(local_pes_23_3_reset),
    .io_in_q(local_pes_23_3_io_in_q),
    .io_in_sum(local_pes_23_3_io_in_sum),
    .io_in_sum_exp(local_pes_23_3_io_in_sum_exp),
    .io_in_kv(local_pes_23_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_3_io_in_inv_sum),
    .io_in_stage(local_pes_23_3_io_in_stage),
    .io_out_q(local_pes_23_3_io_out_q),
    .io_out_sum(local_pes_23_3_io_out_sum),
    .io_out_sum_exp(local_pes_23_3_io_out_sum_exp),
    .io_out_kv(local_pes_23_3_io_out_kv),
    .io_out_stage(local_pes_23_3_io_out_stage)
  );
  PE_1 local_pes_23_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_4_clock),
    .reset(local_pes_23_4_reset),
    .io_in_q(local_pes_23_4_io_in_q),
    .io_in_sum(local_pes_23_4_io_in_sum),
    .io_in_sum_exp(local_pes_23_4_io_in_sum_exp),
    .io_in_kv(local_pes_23_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_4_io_in_inv_sum),
    .io_in_stage(local_pes_23_4_io_in_stage),
    .io_out_q(local_pes_23_4_io_out_q),
    .io_out_sum(local_pes_23_4_io_out_sum),
    .io_out_sum_exp(local_pes_23_4_io_out_sum_exp),
    .io_out_kv(local_pes_23_4_io_out_kv),
    .io_out_stage(local_pes_23_4_io_out_stage)
  );
  PE_1 local_pes_23_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_5_clock),
    .reset(local_pes_23_5_reset),
    .io_in_q(local_pes_23_5_io_in_q),
    .io_in_sum(local_pes_23_5_io_in_sum),
    .io_in_sum_exp(local_pes_23_5_io_in_sum_exp),
    .io_in_kv(local_pes_23_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_5_io_in_inv_sum),
    .io_in_stage(local_pes_23_5_io_in_stage),
    .io_out_q(local_pes_23_5_io_out_q),
    .io_out_sum(local_pes_23_5_io_out_sum),
    .io_out_sum_exp(local_pes_23_5_io_out_sum_exp),
    .io_out_kv(local_pes_23_5_io_out_kv),
    .io_out_stage(local_pes_23_5_io_out_stage)
  );
  PE_1 local_pes_23_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_6_clock),
    .reset(local_pes_23_6_reset),
    .io_in_q(local_pes_23_6_io_in_q),
    .io_in_sum(local_pes_23_6_io_in_sum),
    .io_in_sum_exp(local_pes_23_6_io_in_sum_exp),
    .io_in_kv(local_pes_23_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_6_io_in_inv_sum),
    .io_in_stage(local_pes_23_6_io_in_stage),
    .io_out_q(local_pes_23_6_io_out_q),
    .io_out_sum(local_pes_23_6_io_out_sum),
    .io_out_sum_exp(local_pes_23_6_io_out_sum_exp),
    .io_out_kv(local_pes_23_6_io_out_kv),
    .io_out_stage(local_pes_23_6_io_out_stage)
  );
  PE_1 local_pes_23_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_7_clock),
    .reset(local_pes_23_7_reset),
    .io_in_q(local_pes_23_7_io_in_q),
    .io_in_sum(local_pes_23_7_io_in_sum),
    .io_in_sum_exp(local_pes_23_7_io_in_sum_exp),
    .io_in_kv(local_pes_23_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_7_io_in_inv_sum),
    .io_in_stage(local_pes_23_7_io_in_stage),
    .io_out_q(local_pes_23_7_io_out_q),
    .io_out_sum(local_pes_23_7_io_out_sum),
    .io_out_sum_exp(local_pes_23_7_io_out_sum_exp),
    .io_out_kv(local_pes_23_7_io_out_kv),
    .io_out_stage(local_pes_23_7_io_out_stage)
  );
  PE_1 local_pes_23_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_8_clock),
    .reset(local_pes_23_8_reset),
    .io_in_q(local_pes_23_8_io_in_q),
    .io_in_sum(local_pes_23_8_io_in_sum),
    .io_in_sum_exp(local_pes_23_8_io_in_sum_exp),
    .io_in_kv(local_pes_23_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_8_io_in_inv_sum),
    .io_in_stage(local_pes_23_8_io_in_stage),
    .io_out_q(local_pes_23_8_io_out_q),
    .io_out_sum(local_pes_23_8_io_out_sum),
    .io_out_sum_exp(local_pes_23_8_io_out_sum_exp),
    .io_out_kv(local_pes_23_8_io_out_kv),
    .io_out_stage(local_pes_23_8_io_out_stage)
  );
  PE_1 local_pes_23_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_9_clock),
    .reset(local_pes_23_9_reset),
    .io_in_q(local_pes_23_9_io_in_q),
    .io_in_sum(local_pes_23_9_io_in_sum),
    .io_in_sum_exp(local_pes_23_9_io_in_sum_exp),
    .io_in_kv(local_pes_23_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_9_io_in_inv_sum),
    .io_in_stage(local_pes_23_9_io_in_stage),
    .io_out_q(local_pes_23_9_io_out_q),
    .io_out_sum(local_pes_23_9_io_out_sum),
    .io_out_sum_exp(local_pes_23_9_io_out_sum_exp),
    .io_out_kv(local_pes_23_9_io_out_kv),
    .io_out_stage(local_pes_23_9_io_out_stage)
  );
  PE_1 local_pes_23_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_10_clock),
    .reset(local_pes_23_10_reset),
    .io_in_q(local_pes_23_10_io_in_q),
    .io_in_sum(local_pes_23_10_io_in_sum),
    .io_in_sum_exp(local_pes_23_10_io_in_sum_exp),
    .io_in_kv(local_pes_23_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_10_io_in_inv_sum),
    .io_in_stage(local_pes_23_10_io_in_stage),
    .io_out_q(local_pes_23_10_io_out_q),
    .io_out_sum(local_pes_23_10_io_out_sum),
    .io_out_sum_exp(local_pes_23_10_io_out_sum_exp),
    .io_out_kv(local_pes_23_10_io_out_kv),
    .io_out_stage(local_pes_23_10_io_out_stage)
  );
  PE_1 local_pes_23_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_11_clock),
    .reset(local_pes_23_11_reset),
    .io_in_q(local_pes_23_11_io_in_q),
    .io_in_sum(local_pes_23_11_io_in_sum),
    .io_in_sum_exp(local_pes_23_11_io_in_sum_exp),
    .io_in_kv(local_pes_23_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_11_io_in_inv_sum),
    .io_in_stage(local_pes_23_11_io_in_stage),
    .io_out_q(local_pes_23_11_io_out_q),
    .io_out_sum(local_pes_23_11_io_out_sum),
    .io_out_sum_exp(local_pes_23_11_io_out_sum_exp),
    .io_out_kv(local_pes_23_11_io_out_kv),
    .io_out_stage(local_pes_23_11_io_out_stage)
  );
  PE_1 local_pes_23_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_12_clock),
    .reset(local_pes_23_12_reset),
    .io_in_q(local_pes_23_12_io_in_q),
    .io_in_sum(local_pes_23_12_io_in_sum),
    .io_in_sum_exp(local_pes_23_12_io_in_sum_exp),
    .io_in_kv(local_pes_23_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_12_io_in_inv_sum),
    .io_in_stage(local_pes_23_12_io_in_stage),
    .io_out_q(local_pes_23_12_io_out_q),
    .io_out_sum(local_pes_23_12_io_out_sum),
    .io_out_sum_exp(local_pes_23_12_io_out_sum_exp),
    .io_out_kv(local_pes_23_12_io_out_kv),
    .io_out_stage(local_pes_23_12_io_out_stage)
  );
  PE_1 local_pes_23_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_13_clock),
    .reset(local_pes_23_13_reset),
    .io_in_q(local_pes_23_13_io_in_q),
    .io_in_sum(local_pes_23_13_io_in_sum),
    .io_in_sum_exp(local_pes_23_13_io_in_sum_exp),
    .io_in_kv(local_pes_23_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_13_io_in_inv_sum),
    .io_in_stage(local_pes_23_13_io_in_stage),
    .io_out_q(local_pes_23_13_io_out_q),
    .io_out_sum(local_pes_23_13_io_out_sum),
    .io_out_sum_exp(local_pes_23_13_io_out_sum_exp),
    .io_out_kv(local_pes_23_13_io_out_kv),
    .io_out_stage(local_pes_23_13_io_out_stage)
  );
  PE_1 local_pes_23_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_14_clock),
    .reset(local_pes_23_14_reset),
    .io_in_q(local_pes_23_14_io_in_q),
    .io_in_sum(local_pes_23_14_io_in_sum),
    .io_in_sum_exp(local_pes_23_14_io_in_sum_exp),
    .io_in_kv(local_pes_23_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_14_io_in_inv_sum),
    .io_in_stage(local_pes_23_14_io_in_stage),
    .io_out_q(local_pes_23_14_io_out_q),
    .io_out_sum(local_pes_23_14_io_out_sum),
    .io_out_sum_exp(local_pes_23_14_io_out_sum_exp),
    .io_out_kv(local_pes_23_14_io_out_kv),
    .io_out_stage(local_pes_23_14_io_out_stage)
  );
  PE_1 local_pes_23_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_15_clock),
    .reset(local_pes_23_15_reset),
    .io_in_q(local_pes_23_15_io_in_q),
    .io_in_sum(local_pes_23_15_io_in_sum),
    .io_in_sum_exp(local_pes_23_15_io_in_sum_exp),
    .io_in_kv(local_pes_23_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_15_io_in_inv_sum),
    .io_in_stage(local_pes_23_15_io_in_stage),
    .io_out_q(local_pes_23_15_io_out_q),
    .io_out_sum(local_pes_23_15_io_out_sum),
    .io_out_sum_exp(local_pes_23_15_io_out_sum_exp),
    .io_out_kv(local_pes_23_15_io_out_kv),
    .io_out_stage(local_pes_23_15_io_out_stage)
  );
  PE_1 local_pes_23_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_16_clock),
    .reset(local_pes_23_16_reset),
    .io_in_q(local_pes_23_16_io_in_q),
    .io_in_sum(local_pes_23_16_io_in_sum),
    .io_in_sum_exp(local_pes_23_16_io_in_sum_exp),
    .io_in_kv(local_pes_23_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_16_io_in_inv_sum),
    .io_in_stage(local_pes_23_16_io_in_stage),
    .io_out_q(local_pes_23_16_io_out_q),
    .io_out_sum(local_pes_23_16_io_out_sum),
    .io_out_sum_exp(local_pes_23_16_io_out_sum_exp),
    .io_out_kv(local_pes_23_16_io_out_kv),
    .io_out_stage(local_pes_23_16_io_out_stage)
  );
  PE_1 local_pes_23_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_17_clock),
    .reset(local_pes_23_17_reset),
    .io_in_q(local_pes_23_17_io_in_q),
    .io_in_sum(local_pes_23_17_io_in_sum),
    .io_in_sum_exp(local_pes_23_17_io_in_sum_exp),
    .io_in_kv(local_pes_23_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_17_io_in_inv_sum),
    .io_in_stage(local_pes_23_17_io_in_stage),
    .io_out_q(local_pes_23_17_io_out_q),
    .io_out_sum(local_pes_23_17_io_out_sum),
    .io_out_sum_exp(local_pes_23_17_io_out_sum_exp),
    .io_out_kv(local_pes_23_17_io_out_kv),
    .io_out_stage(local_pes_23_17_io_out_stage)
  );
  PE_1 local_pes_23_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_18_clock),
    .reset(local_pes_23_18_reset),
    .io_in_q(local_pes_23_18_io_in_q),
    .io_in_sum(local_pes_23_18_io_in_sum),
    .io_in_sum_exp(local_pes_23_18_io_in_sum_exp),
    .io_in_kv(local_pes_23_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_18_io_in_inv_sum),
    .io_in_stage(local_pes_23_18_io_in_stage),
    .io_out_q(local_pes_23_18_io_out_q),
    .io_out_sum(local_pes_23_18_io_out_sum),
    .io_out_sum_exp(local_pes_23_18_io_out_sum_exp),
    .io_out_kv(local_pes_23_18_io_out_kv),
    .io_out_stage(local_pes_23_18_io_out_stage)
  );
  PE_1 local_pes_23_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_19_clock),
    .reset(local_pes_23_19_reset),
    .io_in_q(local_pes_23_19_io_in_q),
    .io_in_sum(local_pes_23_19_io_in_sum),
    .io_in_sum_exp(local_pes_23_19_io_in_sum_exp),
    .io_in_kv(local_pes_23_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_19_io_in_inv_sum),
    .io_in_stage(local_pes_23_19_io_in_stage),
    .io_out_q(local_pes_23_19_io_out_q),
    .io_out_sum(local_pes_23_19_io_out_sum),
    .io_out_sum_exp(local_pes_23_19_io_out_sum_exp),
    .io_out_kv(local_pes_23_19_io_out_kv),
    .io_out_stage(local_pes_23_19_io_out_stage)
  );
  PE_1 local_pes_23_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_20_clock),
    .reset(local_pes_23_20_reset),
    .io_in_q(local_pes_23_20_io_in_q),
    .io_in_sum(local_pes_23_20_io_in_sum),
    .io_in_sum_exp(local_pes_23_20_io_in_sum_exp),
    .io_in_kv(local_pes_23_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_20_io_in_inv_sum),
    .io_in_stage(local_pes_23_20_io_in_stage),
    .io_out_q(local_pes_23_20_io_out_q),
    .io_out_sum(local_pes_23_20_io_out_sum),
    .io_out_sum_exp(local_pes_23_20_io_out_sum_exp),
    .io_out_kv(local_pes_23_20_io_out_kv),
    .io_out_stage(local_pes_23_20_io_out_stage)
  );
  PE_1 local_pes_23_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_21_clock),
    .reset(local_pes_23_21_reset),
    .io_in_q(local_pes_23_21_io_in_q),
    .io_in_sum(local_pes_23_21_io_in_sum),
    .io_in_sum_exp(local_pes_23_21_io_in_sum_exp),
    .io_in_kv(local_pes_23_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_21_io_in_inv_sum),
    .io_in_stage(local_pes_23_21_io_in_stage),
    .io_out_q(local_pes_23_21_io_out_q),
    .io_out_sum(local_pes_23_21_io_out_sum),
    .io_out_sum_exp(local_pes_23_21_io_out_sum_exp),
    .io_out_kv(local_pes_23_21_io_out_kv),
    .io_out_stage(local_pes_23_21_io_out_stage)
  );
  PE_1 local_pes_23_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_22_clock),
    .reset(local_pes_23_22_reset),
    .io_in_q(local_pes_23_22_io_in_q),
    .io_in_sum(local_pes_23_22_io_in_sum),
    .io_in_sum_exp(local_pes_23_22_io_in_sum_exp),
    .io_in_kv(local_pes_23_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_22_io_in_inv_sum),
    .io_in_stage(local_pes_23_22_io_in_stage),
    .io_out_q(local_pes_23_22_io_out_q),
    .io_out_sum(local_pes_23_22_io_out_sum),
    .io_out_sum_exp(local_pes_23_22_io_out_sum_exp),
    .io_out_kv(local_pes_23_22_io_out_kv),
    .io_out_stage(local_pes_23_22_io_out_stage)
  );
  PE_1 local_pes_23_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_23_clock),
    .reset(local_pes_23_23_reset),
    .io_in_q(local_pes_23_23_io_in_q),
    .io_in_sum(local_pes_23_23_io_in_sum),
    .io_in_sum_exp(local_pes_23_23_io_in_sum_exp),
    .io_in_kv(local_pes_23_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_23_io_in_inv_sum),
    .io_in_stage(local_pes_23_23_io_in_stage),
    .io_out_q(local_pes_23_23_io_out_q),
    .io_out_sum(local_pes_23_23_io_out_sum),
    .io_out_sum_exp(local_pes_23_23_io_out_sum_exp),
    .io_out_kv(local_pes_23_23_io_out_kv),
    .io_out_stage(local_pes_23_23_io_out_stage)
  );
  PE_1 local_pes_23_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_24_clock),
    .reset(local_pes_23_24_reset),
    .io_in_q(local_pes_23_24_io_in_q),
    .io_in_sum(local_pes_23_24_io_in_sum),
    .io_in_sum_exp(local_pes_23_24_io_in_sum_exp),
    .io_in_kv(local_pes_23_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_24_io_in_inv_sum),
    .io_in_stage(local_pes_23_24_io_in_stage),
    .io_out_q(local_pes_23_24_io_out_q),
    .io_out_sum(local_pes_23_24_io_out_sum),
    .io_out_sum_exp(local_pes_23_24_io_out_sum_exp),
    .io_out_kv(local_pes_23_24_io_out_kv),
    .io_out_stage(local_pes_23_24_io_out_stage)
  );
  PE_1 local_pes_23_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_25_clock),
    .reset(local_pes_23_25_reset),
    .io_in_q(local_pes_23_25_io_in_q),
    .io_in_sum(local_pes_23_25_io_in_sum),
    .io_in_sum_exp(local_pes_23_25_io_in_sum_exp),
    .io_in_kv(local_pes_23_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_25_io_in_inv_sum),
    .io_in_stage(local_pes_23_25_io_in_stage),
    .io_out_q(local_pes_23_25_io_out_q),
    .io_out_sum(local_pes_23_25_io_out_sum),
    .io_out_sum_exp(local_pes_23_25_io_out_sum_exp),
    .io_out_kv(local_pes_23_25_io_out_kv),
    .io_out_stage(local_pes_23_25_io_out_stage)
  );
  PE_1 local_pes_23_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_26_clock),
    .reset(local_pes_23_26_reset),
    .io_in_q(local_pes_23_26_io_in_q),
    .io_in_sum(local_pes_23_26_io_in_sum),
    .io_in_sum_exp(local_pes_23_26_io_in_sum_exp),
    .io_in_kv(local_pes_23_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_26_io_in_inv_sum),
    .io_in_stage(local_pes_23_26_io_in_stage),
    .io_out_q(local_pes_23_26_io_out_q),
    .io_out_sum(local_pes_23_26_io_out_sum),
    .io_out_sum_exp(local_pes_23_26_io_out_sum_exp),
    .io_out_kv(local_pes_23_26_io_out_kv),
    .io_out_stage(local_pes_23_26_io_out_stage)
  );
  PE_1 local_pes_23_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_27_clock),
    .reset(local_pes_23_27_reset),
    .io_in_q(local_pes_23_27_io_in_q),
    .io_in_sum(local_pes_23_27_io_in_sum),
    .io_in_sum_exp(local_pes_23_27_io_in_sum_exp),
    .io_in_kv(local_pes_23_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_27_io_in_inv_sum),
    .io_in_stage(local_pes_23_27_io_in_stage),
    .io_out_q(local_pes_23_27_io_out_q),
    .io_out_sum(local_pes_23_27_io_out_sum),
    .io_out_sum_exp(local_pes_23_27_io_out_sum_exp),
    .io_out_kv(local_pes_23_27_io_out_kv),
    .io_out_stage(local_pes_23_27_io_out_stage)
  );
  PE_1 local_pes_23_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_28_clock),
    .reset(local_pes_23_28_reset),
    .io_in_q(local_pes_23_28_io_in_q),
    .io_in_sum(local_pes_23_28_io_in_sum),
    .io_in_sum_exp(local_pes_23_28_io_in_sum_exp),
    .io_in_kv(local_pes_23_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_28_io_in_inv_sum),
    .io_in_stage(local_pes_23_28_io_in_stage),
    .io_out_q(local_pes_23_28_io_out_q),
    .io_out_sum(local_pes_23_28_io_out_sum),
    .io_out_sum_exp(local_pes_23_28_io_out_sum_exp),
    .io_out_kv(local_pes_23_28_io_out_kv),
    .io_out_stage(local_pes_23_28_io_out_stage)
  );
  PE_1 local_pes_23_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_29_clock),
    .reset(local_pes_23_29_reset),
    .io_in_q(local_pes_23_29_io_in_q),
    .io_in_sum(local_pes_23_29_io_in_sum),
    .io_in_sum_exp(local_pes_23_29_io_in_sum_exp),
    .io_in_kv(local_pes_23_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_29_io_in_inv_sum),
    .io_in_stage(local_pes_23_29_io_in_stage),
    .io_out_q(local_pes_23_29_io_out_q),
    .io_out_sum(local_pes_23_29_io_out_sum),
    .io_out_sum_exp(local_pes_23_29_io_out_sum_exp),
    .io_out_kv(local_pes_23_29_io_out_kv),
    .io_out_stage(local_pes_23_29_io_out_stage)
  );
  PE_1 local_pes_23_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_30_clock),
    .reset(local_pes_23_30_reset),
    .io_in_q(local_pes_23_30_io_in_q),
    .io_in_sum(local_pes_23_30_io_in_sum),
    .io_in_sum_exp(local_pes_23_30_io_in_sum_exp),
    .io_in_kv(local_pes_23_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_30_io_in_inv_sum),
    .io_in_stage(local_pes_23_30_io_in_stage),
    .io_out_q(local_pes_23_30_io_out_q),
    .io_out_sum(local_pes_23_30_io_out_sum),
    .io_out_sum_exp(local_pes_23_30_io_out_sum_exp),
    .io_out_kv(local_pes_23_30_io_out_kv),
    .io_out_stage(local_pes_23_30_io_out_stage)
  );
  PE_1 local_pes_23_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_23_31_clock),
    .reset(local_pes_23_31_reset),
    .io_in_q(local_pes_23_31_io_in_q),
    .io_in_sum(local_pes_23_31_io_in_sum),
    .io_in_sum_exp(local_pes_23_31_io_in_sum_exp),
    .io_in_kv(local_pes_23_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_23_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_23_31_io_in_inv_sum),
    .io_in_stage(local_pes_23_31_io_in_stage),
    .io_out_q(local_pes_23_31_io_out_q),
    .io_out_sum(local_pes_23_31_io_out_sum),
    .io_out_sum_exp(local_pes_23_31_io_out_sum_exp),
    .io_out_kv(local_pes_23_31_io_out_kv),
    .io_out_stage(local_pes_23_31_io_out_stage)
  );
  PE local_pes_24_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_0_clock),
    .reset(local_pes_24_0_reset),
    .io_in_q(local_pes_24_0_io_in_q),
    .io_in_kv(local_pes_24_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_0_io_in_inv_sum),
    .io_in_stage(local_pes_24_0_io_in_stage),
    .io_out_q(local_pes_24_0_io_out_q),
    .io_out_sum(local_pes_24_0_io_out_sum),
    .io_out_kv(local_pes_24_0_io_out_kv),
    .io_out_stage(local_pes_24_0_io_out_stage)
  );
  PE_1 local_pes_24_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_1_clock),
    .reset(local_pes_24_1_reset),
    .io_in_q(local_pes_24_1_io_in_q),
    .io_in_sum(local_pes_24_1_io_in_sum),
    .io_in_sum_exp(local_pes_24_1_io_in_sum_exp),
    .io_in_kv(local_pes_24_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_1_io_in_inv_sum),
    .io_in_stage(local_pes_24_1_io_in_stage),
    .io_out_q(local_pes_24_1_io_out_q),
    .io_out_sum(local_pes_24_1_io_out_sum),
    .io_out_sum_exp(local_pes_24_1_io_out_sum_exp),
    .io_out_kv(local_pes_24_1_io_out_kv),
    .io_out_stage(local_pes_24_1_io_out_stage)
  );
  PE_1 local_pes_24_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_2_clock),
    .reset(local_pes_24_2_reset),
    .io_in_q(local_pes_24_2_io_in_q),
    .io_in_sum(local_pes_24_2_io_in_sum),
    .io_in_sum_exp(local_pes_24_2_io_in_sum_exp),
    .io_in_kv(local_pes_24_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_2_io_in_inv_sum),
    .io_in_stage(local_pes_24_2_io_in_stage),
    .io_out_q(local_pes_24_2_io_out_q),
    .io_out_sum(local_pes_24_2_io_out_sum),
    .io_out_sum_exp(local_pes_24_2_io_out_sum_exp),
    .io_out_kv(local_pes_24_2_io_out_kv),
    .io_out_stage(local_pes_24_2_io_out_stage)
  );
  PE_1 local_pes_24_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_3_clock),
    .reset(local_pes_24_3_reset),
    .io_in_q(local_pes_24_3_io_in_q),
    .io_in_sum(local_pes_24_3_io_in_sum),
    .io_in_sum_exp(local_pes_24_3_io_in_sum_exp),
    .io_in_kv(local_pes_24_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_3_io_in_inv_sum),
    .io_in_stage(local_pes_24_3_io_in_stage),
    .io_out_q(local_pes_24_3_io_out_q),
    .io_out_sum(local_pes_24_3_io_out_sum),
    .io_out_sum_exp(local_pes_24_3_io_out_sum_exp),
    .io_out_kv(local_pes_24_3_io_out_kv),
    .io_out_stage(local_pes_24_3_io_out_stage)
  );
  PE_1 local_pes_24_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_4_clock),
    .reset(local_pes_24_4_reset),
    .io_in_q(local_pes_24_4_io_in_q),
    .io_in_sum(local_pes_24_4_io_in_sum),
    .io_in_sum_exp(local_pes_24_4_io_in_sum_exp),
    .io_in_kv(local_pes_24_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_4_io_in_inv_sum),
    .io_in_stage(local_pes_24_4_io_in_stage),
    .io_out_q(local_pes_24_4_io_out_q),
    .io_out_sum(local_pes_24_4_io_out_sum),
    .io_out_sum_exp(local_pes_24_4_io_out_sum_exp),
    .io_out_kv(local_pes_24_4_io_out_kv),
    .io_out_stage(local_pes_24_4_io_out_stage)
  );
  PE_1 local_pes_24_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_5_clock),
    .reset(local_pes_24_5_reset),
    .io_in_q(local_pes_24_5_io_in_q),
    .io_in_sum(local_pes_24_5_io_in_sum),
    .io_in_sum_exp(local_pes_24_5_io_in_sum_exp),
    .io_in_kv(local_pes_24_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_5_io_in_inv_sum),
    .io_in_stage(local_pes_24_5_io_in_stage),
    .io_out_q(local_pes_24_5_io_out_q),
    .io_out_sum(local_pes_24_5_io_out_sum),
    .io_out_sum_exp(local_pes_24_5_io_out_sum_exp),
    .io_out_kv(local_pes_24_5_io_out_kv),
    .io_out_stage(local_pes_24_5_io_out_stage)
  );
  PE_1 local_pes_24_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_6_clock),
    .reset(local_pes_24_6_reset),
    .io_in_q(local_pes_24_6_io_in_q),
    .io_in_sum(local_pes_24_6_io_in_sum),
    .io_in_sum_exp(local_pes_24_6_io_in_sum_exp),
    .io_in_kv(local_pes_24_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_6_io_in_inv_sum),
    .io_in_stage(local_pes_24_6_io_in_stage),
    .io_out_q(local_pes_24_6_io_out_q),
    .io_out_sum(local_pes_24_6_io_out_sum),
    .io_out_sum_exp(local_pes_24_6_io_out_sum_exp),
    .io_out_kv(local_pes_24_6_io_out_kv),
    .io_out_stage(local_pes_24_6_io_out_stage)
  );
  PE_1 local_pes_24_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_7_clock),
    .reset(local_pes_24_7_reset),
    .io_in_q(local_pes_24_7_io_in_q),
    .io_in_sum(local_pes_24_7_io_in_sum),
    .io_in_sum_exp(local_pes_24_7_io_in_sum_exp),
    .io_in_kv(local_pes_24_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_7_io_in_inv_sum),
    .io_in_stage(local_pes_24_7_io_in_stage),
    .io_out_q(local_pes_24_7_io_out_q),
    .io_out_sum(local_pes_24_7_io_out_sum),
    .io_out_sum_exp(local_pes_24_7_io_out_sum_exp),
    .io_out_kv(local_pes_24_7_io_out_kv),
    .io_out_stage(local_pes_24_7_io_out_stage)
  );
  PE_1 local_pes_24_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_8_clock),
    .reset(local_pes_24_8_reset),
    .io_in_q(local_pes_24_8_io_in_q),
    .io_in_sum(local_pes_24_8_io_in_sum),
    .io_in_sum_exp(local_pes_24_8_io_in_sum_exp),
    .io_in_kv(local_pes_24_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_8_io_in_inv_sum),
    .io_in_stage(local_pes_24_8_io_in_stage),
    .io_out_q(local_pes_24_8_io_out_q),
    .io_out_sum(local_pes_24_8_io_out_sum),
    .io_out_sum_exp(local_pes_24_8_io_out_sum_exp),
    .io_out_kv(local_pes_24_8_io_out_kv),
    .io_out_stage(local_pes_24_8_io_out_stage)
  );
  PE_1 local_pes_24_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_9_clock),
    .reset(local_pes_24_9_reset),
    .io_in_q(local_pes_24_9_io_in_q),
    .io_in_sum(local_pes_24_9_io_in_sum),
    .io_in_sum_exp(local_pes_24_9_io_in_sum_exp),
    .io_in_kv(local_pes_24_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_9_io_in_inv_sum),
    .io_in_stage(local_pes_24_9_io_in_stage),
    .io_out_q(local_pes_24_9_io_out_q),
    .io_out_sum(local_pes_24_9_io_out_sum),
    .io_out_sum_exp(local_pes_24_9_io_out_sum_exp),
    .io_out_kv(local_pes_24_9_io_out_kv),
    .io_out_stage(local_pes_24_9_io_out_stage)
  );
  PE_1 local_pes_24_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_10_clock),
    .reset(local_pes_24_10_reset),
    .io_in_q(local_pes_24_10_io_in_q),
    .io_in_sum(local_pes_24_10_io_in_sum),
    .io_in_sum_exp(local_pes_24_10_io_in_sum_exp),
    .io_in_kv(local_pes_24_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_10_io_in_inv_sum),
    .io_in_stage(local_pes_24_10_io_in_stage),
    .io_out_q(local_pes_24_10_io_out_q),
    .io_out_sum(local_pes_24_10_io_out_sum),
    .io_out_sum_exp(local_pes_24_10_io_out_sum_exp),
    .io_out_kv(local_pes_24_10_io_out_kv),
    .io_out_stage(local_pes_24_10_io_out_stage)
  );
  PE_1 local_pes_24_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_11_clock),
    .reset(local_pes_24_11_reset),
    .io_in_q(local_pes_24_11_io_in_q),
    .io_in_sum(local_pes_24_11_io_in_sum),
    .io_in_sum_exp(local_pes_24_11_io_in_sum_exp),
    .io_in_kv(local_pes_24_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_11_io_in_inv_sum),
    .io_in_stage(local_pes_24_11_io_in_stage),
    .io_out_q(local_pes_24_11_io_out_q),
    .io_out_sum(local_pes_24_11_io_out_sum),
    .io_out_sum_exp(local_pes_24_11_io_out_sum_exp),
    .io_out_kv(local_pes_24_11_io_out_kv),
    .io_out_stage(local_pes_24_11_io_out_stage)
  );
  PE_1 local_pes_24_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_12_clock),
    .reset(local_pes_24_12_reset),
    .io_in_q(local_pes_24_12_io_in_q),
    .io_in_sum(local_pes_24_12_io_in_sum),
    .io_in_sum_exp(local_pes_24_12_io_in_sum_exp),
    .io_in_kv(local_pes_24_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_12_io_in_inv_sum),
    .io_in_stage(local_pes_24_12_io_in_stage),
    .io_out_q(local_pes_24_12_io_out_q),
    .io_out_sum(local_pes_24_12_io_out_sum),
    .io_out_sum_exp(local_pes_24_12_io_out_sum_exp),
    .io_out_kv(local_pes_24_12_io_out_kv),
    .io_out_stage(local_pes_24_12_io_out_stage)
  );
  PE_1 local_pes_24_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_13_clock),
    .reset(local_pes_24_13_reset),
    .io_in_q(local_pes_24_13_io_in_q),
    .io_in_sum(local_pes_24_13_io_in_sum),
    .io_in_sum_exp(local_pes_24_13_io_in_sum_exp),
    .io_in_kv(local_pes_24_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_13_io_in_inv_sum),
    .io_in_stage(local_pes_24_13_io_in_stage),
    .io_out_q(local_pes_24_13_io_out_q),
    .io_out_sum(local_pes_24_13_io_out_sum),
    .io_out_sum_exp(local_pes_24_13_io_out_sum_exp),
    .io_out_kv(local_pes_24_13_io_out_kv),
    .io_out_stage(local_pes_24_13_io_out_stage)
  );
  PE_1 local_pes_24_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_14_clock),
    .reset(local_pes_24_14_reset),
    .io_in_q(local_pes_24_14_io_in_q),
    .io_in_sum(local_pes_24_14_io_in_sum),
    .io_in_sum_exp(local_pes_24_14_io_in_sum_exp),
    .io_in_kv(local_pes_24_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_14_io_in_inv_sum),
    .io_in_stage(local_pes_24_14_io_in_stage),
    .io_out_q(local_pes_24_14_io_out_q),
    .io_out_sum(local_pes_24_14_io_out_sum),
    .io_out_sum_exp(local_pes_24_14_io_out_sum_exp),
    .io_out_kv(local_pes_24_14_io_out_kv),
    .io_out_stage(local_pes_24_14_io_out_stage)
  );
  PE_1 local_pes_24_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_15_clock),
    .reset(local_pes_24_15_reset),
    .io_in_q(local_pes_24_15_io_in_q),
    .io_in_sum(local_pes_24_15_io_in_sum),
    .io_in_sum_exp(local_pes_24_15_io_in_sum_exp),
    .io_in_kv(local_pes_24_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_15_io_in_inv_sum),
    .io_in_stage(local_pes_24_15_io_in_stage),
    .io_out_q(local_pes_24_15_io_out_q),
    .io_out_sum(local_pes_24_15_io_out_sum),
    .io_out_sum_exp(local_pes_24_15_io_out_sum_exp),
    .io_out_kv(local_pes_24_15_io_out_kv),
    .io_out_stage(local_pes_24_15_io_out_stage)
  );
  PE_1 local_pes_24_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_16_clock),
    .reset(local_pes_24_16_reset),
    .io_in_q(local_pes_24_16_io_in_q),
    .io_in_sum(local_pes_24_16_io_in_sum),
    .io_in_sum_exp(local_pes_24_16_io_in_sum_exp),
    .io_in_kv(local_pes_24_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_16_io_in_inv_sum),
    .io_in_stage(local_pes_24_16_io_in_stage),
    .io_out_q(local_pes_24_16_io_out_q),
    .io_out_sum(local_pes_24_16_io_out_sum),
    .io_out_sum_exp(local_pes_24_16_io_out_sum_exp),
    .io_out_kv(local_pes_24_16_io_out_kv),
    .io_out_stage(local_pes_24_16_io_out_stage)
  );
  PE_1 local_pes_24_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_17_clock),
    .reset(local_pes_24_17_reset),
    .io_in_q(local_pes_24_17_io_in_q),
    .io_in_sum(local_pes_24_17_io_in_sum),
    .io_in_sum_exp(local_pes_24_17_io_in_sum_exp),
    .io_in_kv(local_pes_24_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_17_io_in_inv_sum),
    .io_in_stage(local_pes_24_17_io_in_stage),
    .io_out_q(local_pes_24_17_io_out_q),
    .io_out_sum(local_pes_24_17_io_out_sum),
    .io_out_sum_exp(local_pes_24_17_io_out_sum_exp),
    .io_out_kv(local_pes_24_17_io_out_kv),
    .io_out_stage(local_pes_24_17_io_out_stage)
  );
  PE_1 local_pes_24_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_18_clock),
    .reset(local_pes_24_18_reset),
    .io_in_q(local_pes_24_18_io_in_q),
    .io_in_sum(local_pes_24_18_io_in_sum),
    .io_in_sum_exp(local_pes_24_18_io_in_sum_exp),
    .io_in_kv(local_pes_24_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_18_io_in_inv_sum),
    .io_in_stage(local_pes_24_18_io_in_stage),
    .io_out_q(local_pes_24_18_io_out_q),
    .io_out_sum(local_pes_24_18_io_out_sum),
    .io_out_sum_exp(local_pes_24_18_io_out_sum_exp),
    .io_out_kv(local_pes_24_18_io_out_kv),
    .io_out_stage(local_pes_24_18_io_out_stage)
  );
  PE_1 local_pes_24_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_19_clock),
    .reset(local_pes_24_19_reset),
    .io_in_q(local_pes_24_19_io_in_q),
    .io_in_sum(local_pes_24_19_io_in_sum),
    .io_in_sum_exp(local_pes_24_19_io_in_sum_exp),
    .io_in_kv(local_pes_24_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_19_io_in_inv_sum),
    .io_in_stage(local_pes_24_19_io_in_stage),
    .io_out_q(local_pes_24_19_io_out_q),
    .io_out_sum(local_pes_24_19_io_out_sum),
    .io_out_sum_exp(local_pes_24_19_io_out_sum_exp),
    .io_out_kv(local_pes_24_19_io_out_kv),
    .io_out_stage(local_pes_24_19_io_out_stage)
  );
  PE_1 local_pes_24_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_20_clock),
    .reset(local_pes_24_20_reset),
    .io_in_q(local_pes_24_20_io_in_q),
    .io_in_sum(local_pes_24_20_io_in_sum),
    .io_in_sum_exp(local_pes_24_20_io_in_sum_exp),
    .io_in_kv(local_pes_24_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_20_io_in_inv_sum),
    .io_in_stage(local_pes_24_20_io_in_stage),
    .io_out_q(local_pes_24_20_io_out_q),
    .io_out_sum(local_pes_24_20_io_out_sum),
    .io_out_sum_exp(local_pes_24_20_io_out_sum_exp),
    .io_out_kv(local_pes_24_20_io_out_kv),
    .io_out_stage(local_pes_24_20_io_out_stage)
  );
  PE_1 local_pes_24_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_21_clock),
    .reset(local_pes_24_21_reset),
    .io_in_q(local_pes_24_21_io_in_q),
    .io_in_sum(local_pes_24_21_io_in_sum),
    .io_in_sum_exp(local_pes_24_21_io_in_sum_exp),
    .io_in_kv(local_pes_24_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_21_io_in_inv_sum),
    .io_in_stage(local_pes_24_21_io_in_stage),
    .io_out_q(local_pes_24_21_io_out_q),
    .io_out_sum(local_pes_24_21_io_out_sum),
    .io_out_sum_exp(local_pes_24_21_io_out_sum_exp),
    .io_out_kv(local_pes_24_21_io_out_kv),
    .io_out_stage(local_pes_24_21_io_out_stage)
  );
  PE_1 local_pes_24_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_22_clock),
    .reset(local_pes_24_22_reset),
    .io_in_q(local_pes_24_22_io_in_q),
    .io_in_sum(local_pes_24_22_io_in_sum),
    .io_in_sum_exp(local_pes_24_22_io_in_sum_exp),
    .io_in_kv(local_pes_24_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_22_io_in_inv_sum),
    .io_in_stage(local_pes_24_22_io_in_stage),
    .io_out_q(local_pes_24_22_io_out_q),
    .io_out_sum(local_pes_24_22_io_out_sum),
    .io_out_sum_exp(local_pes_24_22_io_out_sum_exp),
    .io_out_kv(local_pes_24_22_io_out_kv),
    .io_out_stage(local_pes_24_22_io_out_stage)
  );
  PE_1 local_pes_24_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_23_clock),
    .reset(local_pes_24_23_reset),
    .io_in_q(local_pes_24_23_io_in_q),
    .io_in_sum(local_pes_24_23_io_in_sum),
    .io_in_sum_exp(local_pes_24_23_io_in_sum_exp),
    .io_in_kv(local_pes_24_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_23_io_in_inv_sum),
    .io_in_stage(local_pes_24_23_io_in_stage),
    .io_out_q(local_pes_24_23_io_out_q),
    .io_out_sum(local_pes_24_23_io_out_sum),
    .io_out_sum_exp(local_pes_24_23_io_out_sum_exp),
    .io_out_kv(local_pes_24_23_io_out_kv),
    .io_out_stage(local_pes_24_23_io_out_stage)
  );
  PE_1 local_pes_24_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_24_clock),
    .reset(local_pes_24_24_reset),
    .io_in_q(local_pes_24_24_io_in_q),
    .io_in_sum(local_pes_24_24_io_in_sum),
    .io_in_sum_exp(local_pes_24_24_io_in_sum_exp),
    .io_in_kv(local_pes_24_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_24_io_in_inv_sum),
    .io_in_stage(local_pes_24_24_io_in_stage),
    .io_out_q(local_pes_24_24_io_out_q),
    .io_out_sum(local_pes_24_24_io_out_sum),
    .io_out_sum_exp(local_pes_24_24_io_out_sum_exp),
    .io_out_kv(local_pes_24_24_io_out_kv),
    .io_out_stage(local_pes_24_24_io_out_stage)
  );
  PE_1 local_pes_24_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_25_clock),
    .reset(local_pes_24_25_reset),
    .io_in_q(local_pes_24_25_io_in_q),
    .io_in_sum(local_pes_24_25_io_in_sum),
    .io_in_sum_exp(local_pes_24_25_io_in_sum_exp),
    .io_in_kv(local_pes_24_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_25_io_in_inv_sum),
    .io_in_stage(local_pes_24_25_io_in_stage),
    .io_out_q(local_pes_24_25_io_out_q),
    .io_out_sum(local_pes_24_25_io_out_sum),
    .io_out_sum_exp(local_pes_24_25_io_out_sum_exp),
    .io_out_kv(local_pes_24_25_io_out_kv),
    .io_out_stage(local_pes_24_25_io_out_stage)
  );
  PE_1 local_pes_24_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_26_clock),
    .reset(local_pes_24_26_reset),
    .io_in_q(local_pes_24_26_io_in_q),
    .io_in_sum(local_pes_24_26_io_in_sum),
    .io_in_sum_exp(local_pes_24_26_io_in_sum_exp),
    .io_in_kv(local_pes_24_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_26_io_in_inv_sum),
    .io_in_stage(local_pes_24_26_io_in_stage),
    .io_out_q(local_pes_24_26_io_out_q),
    .io_out_sum(local_pes_24_26_io_out_sum),
    .io_out_sum_exp(local_pes_24_26_io_out_sum_exp),
    .io_out_kv(local_pes_24_26_io_out_kv),
    .io_out_stage(local_pes_24_26_io_out_stage)
  );
  PE_1 local_pes_24_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_27_clock),
    .reset(local_pes_24_27_reset),
    .io_in_q(local_pes_24_27_io_in_q),
    .io_in_sum(local_pes_24_27_io_in_sum),
    .io_in_sum_exp(local_pes_24_27_io_in_sum_exp),
    .io_in_kv(local_pes_24_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_27_io_in_inv_sum),
    .io_in_stage(local_pes_24_27_io_in_stage),
    .io_out_q(local_pes_24_27_io_out_q),
    .io_out_sum(local_pes_24_27_io_out_sum),
    .io_out_sum_exp(local_pes_24_27_io_out_sum_exp),
    .io_out_kv(local_pes_24_27_io_out_kv),
    .io_out_stage(local_pes_24_27_io_out_stage)
  );
  PE_1 local_pes_24_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_28_clock),
    .reset(local_pes_24_28_reset),
    .io_in_q(local_pes_24_28_io_in_q),
    .io_in_sum(local_pes_24_28_io_in_sum),
    .io_in_sum_exp(local_pes_24_28_io_in_sum_exp),
    .io_in_kv(local_pes_24_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_28_io_in_inv_sum),
    .io_in_stage(local_pes_24_28_io_in_stage),
    .io_out_q(local_pes_24_28_io_out_q),
    .io_out_sum(local_pes_24_28_io_out_sum),
    .io_out_sum_exp(local_pes_24_28_io_out_sum_exp),
    .io_out_kv(local_pes_24_28_io_out_kv),
    .io_out_stage(local_pes_24_28_io_out_stage)
  );
  PE_1 local_pes_24_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_29_clock),
    .reset(local_pes_24_29_reset),
    .io_in_q(local_pes_24_29_io_in_q),
    .io_in_sum(local_pes_24_29_io_in_sum),
    .io_in_sum_exp(local_pes_24_29_io_in_sum_exp),
    .io_in_kv(local_pes_24_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_29_io_in_inv_sum),
    .io_in_stage(local_pes_24_29_io_in_stage),
    .io_out_q(local_pes_24_29_io_out_q),
    .io_out_sum(local_pes_24_29_io_out_sum),
    .io_out_sum_exp(local_pes_24_29_io_out_sum_exp),
    .io_out_kv(local_pes_24_29_io_out_kv),
    .io_out_stage(local_pes_24_29_io_out_stage)
  );
  PE_1 local_pes_24_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_30_clock),
    .reset(local_pes_24_30_reset),
    .io_in_q(local_pes_24_30_io_in_q),
    .io_in_sum(local_pes_24_30_io_in_sum),
    .io_in_sum_exp(local_pes_24_30_io_in_sum_exp),
    .io_in_kv(local_pes_24_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_30_io_in_inv_sum),
    .io_in_stage(local_pes_24_30_io_in_stage),
    .io_out_q(local_pes_24_30_io_out_q),
    .io_out_sum(local_pes_24_30_io_out_sum),
    .io_out_sum_exp(local_pes_24_30_io_out_sum_exp),
    .io_out_kv(local_pes_24_30_io_out_kv),
    .io_out_stage(local_pes_24_30_io_out_stage)
  );
  PE_1 local_pes_24_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_24_31_clock),
    .reset(local_pes_24_31_reset),
    .io_in_q(local_pes_24_31_io_in_q),
    .io_in_sum(local_pes_24_31_io_in_sum),
    .io_in_sum_exp(local_pes_24_31_io_in_sum_exp),
    .io_in_kv(local_pes_24_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_24_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_24_31_io_in_inv_sum),
    .io_in_stage(local_pes_24_31_io_in_stage),
    .io_out_q(local_pes_24_31_io_out_q),
    .io_out_sum(local_pes_24_31_io_out_sum),
    .io_out_sum_exp(local_pes_24_31_io_out_sum_exp),
    .io_out_kv(local_pes_24_31_io_out_kv),
    .io_out_stage(local_pes_24_31_io_out_stage)
  );
  PE local_pes_25_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_0_clock),
    .reset(local_pes_25_0_reset),
    .io_in_q(local_pes_25_0_io_in_q),
    .io_in_kv(local_pes_25_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_0_io_in_inv_sum),
    .io_in_stage(local_pes_25_0_io_in_stage),
    .io_out_q(local_pes_25_0_io_out_q),
    .io_out_sum(local_pes_25_0_io_out_sum),
    .io_out_kv(local_pes_25_0_io_out_kv),
    .io_out_stage(local_pes_25_0_io_out_stage)
  );
  PE_1 local_pes_25_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_1_clock),
    .reset(local_pes_25_1_reset),
    .io_in_q(local_pes_25_1_io_in_q),
    .io_in_sum(local_pes_25_1_io_in_sum),
    .io_in_sum_exp(local_pes_25_1_io_in_sum_exp),
    .io_in_kv(local_pes_25_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_1_io_in_inv_sum),
    .io_in_stage(local_pes_25_1_io_in_stage),
    .io_out_q(local_pes_25_1_io_out_q),
    .io_out_sum(local_pes_25_1_io_out_sum),
    .io_out_sum_exp(local_pes_25_1_io_out_sum_exp),
    .io_out_kv(local_pes_25_1_io_out_kv),
    .io_out_stage(local_pes_25_1_io_out_stage)
  );
  PE_1 local_pes_25_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_2_clock),
    .reset(local_pes_25_2_reset),
    .io_in_q(local_pes_25_2_io_in_q),
    .io_in_sum(local_pes_25_2_io_in_sum),
    .io_in_sum_exp(local_pes_25_2_io_in_sum_exp),
    .io_in_kv(local_pes_25_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_2_io_in_inv_sum),
    .io_in_stage(local_pes_25_2_io_in_stage),
    .io_out_q(local_pes_25_2_io_out_q),
    .io_out_sum(local_pes_25_2_io_out_sum),
    .io_out_sum_exp(local_pes_25_2_io_out_sum_exp),
    .io_out_kv(local_pes_25_2_io_out_kv),
    .io_out_stage(local_pes_25_2_io_out_stage)
  );
  PE_1 local_pes_25_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_3_clock),
    .reset(local_pes_25_3_reset),
    .io_in_q(local_pes_25_3_io_in_q),
    .io_in_sum(local_pes_25_3_io_in_sum),
    .io_in_sum_exp(local_pes_25_3_io_in_sum_exp),
    .io_in_kv(local_pes_25_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_3_io_in_inv_sum),
    .io_in_stage(local_pes_25_3_io_in_stage),
    .io_out_q(local_pes_25_3_io_out_q),
    .io_out_sum(local_pes_25_3_io_out_sum),
    .io_out_sum_exp(local_pes_25_3_io_out_sum_exp),
    .io_out_kv(local_pes_25_3_io_out_kv),
    .io_out_stage(local_pes_25_3_io_out_stage)
  );
  PE_1 local_pes_25_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_4_clock),
    .reset(local_pes_25_4_reset),
    .io_in_q(local_pes_25_4_io_in_q),
    .io_in_sum(local_pes_25_4_io_in_sum),
    .io_in_sum_exp(local_pes_25_4_io_in_sum_exp),
    .io_in_kv(local_pes_25_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_4_io_in_inv_sum),
    .io_in_stage(local_pes_25_4_io_in_stage),
    .io_out_q(local_pes_25_4_io_out_q),
    .io_out_sum(local_pes_25_4_io_out_sum),
    .io_out_sum_exp(local_pes_25_4_io_out_sum_exp),
    .io_out_kv(local_pes_25_4_io_out_kv),
    .io_out_stage(local_pes_25_4_io_out_stage)
  );
  PE_1 local_pes_25_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_5_clock),
    .reset(local_pes_25_5_reset),
    .io_in_q(local_pes_25_5_io_in_q),
    .io_in_sum(local_pes_25_5_io_in_sum),
    .io_in_sum_exp(local_pes_25_5_io_in_sum_exp),
    .io_in_kv(local_pes_25_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_5_io_in_inv_sum),
    .io_in_stage(local_pes_25_5_io_in_stage),
    .io_out_q(local_pes_25_5_io_out_q),
    .io_out_sum(local_pes_25_5_io_out_sum),
    .io_out_sum_exp(local_pes_25_5_io_out_sum_exp),
    .io_out_kv(local_pes_25_5_io_out_kv),
    .io_out_stage(local_pes_25_5_io_out_stage)
  );
  PE_1 local_pes_25_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_6_clock),
    .reset(local_pes_25_6_reset),
    .io_in_q(local_pes_25_6_io_in_q),
    .io_in_sum(local_pes_25_6_io_in_sum),
    .io_in_sum_exp(local_pes_25_6_io_in_sum_exp),
    .io_in_kv(local_pes_25_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_6_io_in_inv_sum),
    .io_in_stage(local_pes_25_6_io_in_stage),
    .io_out_q(local_pes_25_6_io_out_q),
    .io_out_sum(local_pes_25_6_io_out_sum),
    .io_out_sum_exp(local_pes_25_6_io_out_sum_exp),
    .io_out_kv(local_pes_25_6_io_out_kv),
    .io_out_stage(local_pes_25_6_io_out_stage)
  );
  PE_1 local_pes_25_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_7_clock),
    .reset(local_pes_25_7_reset),
    .io_in_q(local_pes_25_7_io_in_q),
    .io_in_sum(local_pes_25_7_io_in_sum),
    .io_in_sum_exp(local_pes_25_7_io_in_sum_exp),
    .io_in_kv(local_pes_25_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_7_io_in_inv_sum),
    .io_in_stage(local_pes_25_7_io_in_stage),
    .io_out_q(local_pes_25_7_io_out_q),
    .io_out_sum(local_pes_25_7_io_out_sum),
    .io_out_sum_exp(local_pes_25_7_io_out_sum_exp),
    .io_out_kv(local_pes_25_7_io_out_kv),
    .io_out_stage(local_pes_25_7_io_out_stage)
  );
  PE_1 local_pes_25_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_8_clock),
    .reset(local_pes_25_8_reset),
    .io_in_q(local_pes_25_8_io_in_q),
    .io_in_sum(local_pes_25_8_io_in_sum),
    .io_in_sum_exp(local_pes_25_8_io_in_sum_exp),
    .io_in_kv(local_pes_25_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_8_io_in_inv_sum),
    .io_in_stage(local_pes_25_8_io_in_stage),
    .io_out_q(local_pes_25_8_io_out_q),
    .io_out_sum(local_pes_25_8_io_out_sum),
    .io_out_sum_exp(local_pes_25_8_io_out_sum_exp),
    .io_out_kv(local_pes_25_8_io_out_kv),
    .io_out_stage(local_pes_25_8_io_out_stage)
  );
  PE_1 local_pes_25_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_9_clock),
    .reset(local_pes_25_9_reset),
    .io_in_q(local_pes_25_9_io_in_q),
    .io_in_sum(local_pes_25_9_io_in_sum),
    .io_in_sum_exp(local_pes_25_9_io_in_sum_exp),
    .io_in_kv(local_pes_25_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_9_io_in_inv_sum),
    .io_in_stage(local_pes_25_9_io_in_stage),
    .io_out_q(local_pes_25_9_io_out_q),
    .io_out_sum(local_pes_25_9_io_out_sum),
    .io_out_sum_exp(local_pes_25_9_io_out_sum_exp),
    .io_out_kv(local_pes_25_9_io_out_kv),
    .io_out_stage(local_pes_25_9_io_out_stage)
  );
  PE_1 local_pes_25_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_10_clock),
    .reset(local_pes_25_10_reset),
    .io_in_q(local_pes_25_10_io_in_q),
    .io_in_sum(local_pes_25_10_io_in_sum),
    .io_in_sum_exp(local_pes_25_10_io_in_sum_exp),
    .io_in_kv(local_pes_25_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_10_io_in_inv_sum),
    .io_in_stage(local_pes_25_10_io_in_stage),
    .io_out_q(local_pes_25_10_io_out_q),
    .io_out_sum(local_pes_25_10_io_out_sum),
    .io_out_sum_exp(local_pes_25_10_io_out_sum_exp),
    .io_out_kv(local_pes_25_10_io_out_kv),
    .io_out_stage(local_pes_25_10_io_out_stage)
  );
  PE_1 local_pes_25_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_11_clock),
    .reset(local_pes_25_11_reset),
    .io_in_q(local_pes_25_11_io_in_q),
    .io_in_sum(local_pes_25_11_io_in_sum),
    .io_in_sum_exp(local_pes_25_11_io_in_sum_exp),
    .io_in_kv(local_pes_25_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_11_io_in_inv_sum),
    .io_in_stage(local_pes_25_11_io_in_stage),
    .io_out_q(local_pes_25_11_io_out_q),
    .io_out_sum(local_pes_25_11_io_out_sum),
    .io_out_sum_exp(local_pes_25_11_io_out_sum_exp),
    .io_out_kv(local_pes_25_11_io_out_kv),
    .io_out_stage(local_pes_25_11_io_out_stage)
  );
  PE_1 local_pes_25_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_12_clock),
    .reset(local_pes_25_12_reset),
    .io_in_q(local_pes_25_12_io_in_q),
    .io_in_sum(local_pes_25_12_io_in_sum),
    .io_in_sum_exp(local_pes_25_12_io_in_sum_exp),
    .io_in_kv(local_pes_25_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_12_io_in_inv_sum),
    .io_in_stage(local_pes_25_12_io_in_stage),
    .io_out_q(local_pes_25_12_io_out_q),
    .io_out_sum(local_pes_25_12_io_out_sum),
    .io_out_sum_exp(local_pes_25_12_io_out_sum_exp),
    .io_out_kv(local_pes_25_12_io_out_kv),
    .io_out_stage(local_pes_25_12_io_out_stage)
  );
  PE_1 local_pes_25_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_13_clock),
    .reset(local_pes_25_13_reset),
    .io_in_q(local_pes_25_13_io_in_q),
    .io_in_sum(local_pes_25_13_io_in_sum),
    .io_in_sum_exp(local_pes_25_13_io_in_sum_exp),
    .io_in_kv(local_pes_25_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_13_io_in_inv_sum),
    .io_in_stage(local_pes_25_13_io_in_stage),
    .io_out_q(local_pes_25_13_io_out_q),
    .io_out_sum(local_pes_25_13_io_out_sum),
    .io_out_sum_exp(local_pes_25_13_io_out_sum_exp),
    .io_out_kv(local_pes_25_13_io_out_kv),
    .io_out_stage(local_pes_25_13_io_out_stage)
  );
  PE_1 local_pes_25_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_14_clock),
    .reset(local_pes_25_14_reset),
    .io_in_q(local_pes_25_14_io_in_q),
    .io_in_sum(local_pes_25_14_io_in_sum),
    .io_in_sum_exp(local_pes_25_14_io_in_sum_exp),
    .io_in_kv(local_pes_25_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_14_io_in_inv_sum),
    .io_in_stage(local_pes_25_14_io_in_stage),
    .io_out_q(local_pes_25_14_io_out_q),
    .io_out_sum(local_pes_25_14_io_out_sum),
    .io_out_sum_exp(local_pes_25_14_io_out_sum_exp),
    .io_out_kv(local_pes_25_14_io_out_kv),
    .io_out_stage(local_pes_25_14_io_out_stage)
  );
  PE_1 local_pes_25_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_15_clock),
    .reset(local_pes_25_15_reset),
    .io_in_q(local_pes_25_15_io_in_q),
    .io_in_sum(local_pes_25_15_io_in_sum),
    .io_in_sum_exp(local_pes_25_15_io_in_sum_exp),
    .io_in_kv(local_pes_25_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_15_io_in_inv_sum),
    .io_in_stage(local_pes_25_15_io_in_stage),
    .io_out_q(local_pes_25_15_io_out_q),
    .io_out_sum(local_pes_25_15_io_out_sum),
    .io_out_sum_exp(local_pes_25_15_io_out_sum_exp),
    .io_out_kv(local_pes_25_15_io_out_kv),
    .io_out_stage(local_pes_25_15_io_out_stage)
  );
  PE_1 local_pes_25_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_16_clock),
    .reset(local_pes_25_16_reset),
    .io_in_q(local_pes_25_16_io_in_q),
    .io_in_sum(local_pes_25_16_io_in_sum),
    .io_in_sum_exp(local_pes_25_16_io_in_sum_exp),
    .io_in_kv(local_pes_25_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_16_io_in_inv_sum),
    .io_in_stage(local_pes_25_16_io_in_stage),
    .io_out_q(local_pes_25_16_io_out_q),
    .io_out_sum(local_pes_25_16_io_out_sum),
    .io_out_sum_exp(local_pes_25_16_io_out_sum_exp),
    .io_out_kv(local_pes_25_16_io_out_kv),
    .io_out_stage(local_pes_25_16_io_out_stage)
  );
  PE_1 local_pes_25_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_17_clock),
    .reset(local_pes_25_17_reset),
    .io_in_q(local_pes_25_17_io_in_q),
    .io_in_sum(local_pes_25_17_io_in_sum),
    .io_in_sum_exp(local_pes_25_17_io_in_sum_exp),
    .io_in_kv(local_pes_25_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_17_io_in_inv_sum),
    .io_in_stage(local_pes_25_17_io_in_stage),
    .io_out_q(local_pes_25_17_io_out_q),
    .io_out_sum(local_pes_25_17_io_out_sum),
    .io_out_sum_exp(local_pes_25_17_io_out_sum_exp),
    .io_out_kv(local_pes_25_17_io_out_kv),
    .io_out_stage(local_pes_25_17_io_out_stage)
  );
  PE_1 local_pes_25_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_18_clock),
    .reset(local_pes_25_18_reset),
    .io_in_q(local_pes_25_18_io_in_q),
    .io_in_sum(local_pes_25_18_io_in_sum),
    .io_in_sum_exp(local_pes_25_18_io_in_sum_exp),
    .io_in_kv(local_pes_25_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_18_io_in_inv_sum),
    .io_in_stage(local_pes_25_18_io_in_stage),
    .io_out_q(local_pes_25_18_io_out_q),
    .io_out_sum(local_pes_25_18_io_out_sum),
    .io_out_sum_exp(local_pes_25_18_io_out_sum_exp),
    .io_out_kv(local_pes_25_18_io_out_kv),
    .io_out_stage(local_pes_25_18_io_out_stage)
  );
  PE_1 local_pes_25_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_19_clock),
    .reset(local_pes_25_19_reset),
    .io_in_q(local_pes_25_19_io_in_q),
    .io_in_sum(local_pes_25_19_io_in_sum),
    .io_in_sum_exp(local_pes_25_19_io_in_sum_exp),
    .io_in_kv(local_pes_25_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_19_io_in_inv_sum),
    .io_in_stage(local_pes_25_19_io_in_stage),
    .io_out_q(local_pes_25_19_io_out_q),
    .io_out_sum(local_pes_25_19_io_out_sum),
    .io_out_sum_exp(local_pes_25_19_io_out_sum_exp),
    .io_out_kv(local_pes_25_19_io_out_kv),
    .io_out_stage(local_pes_25_19_io_out_stage)
  );
  PE_1 local_pes_25_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_20_clock),
    .reset(local_pes_25_20_reset),
    .io_in_q(local_pes_25_20_io_in_q),
    .io_in_sum(local_pes_25_20_io_in_sum),
    .io_in_sum_exp(local_pes_25_20_io_in_sum_exp),
    .io_in_kv(local_pes_25_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_20_io_in_inv_sum),
    .io_in_stage(local_pes_25_20_io_in_stage),
    .io_out_q(local_pes_25_20_io_out_q),
    .io_out_sum(local_pes_25_20_io_out_sum),
    .io_out_sum_exp(local_pes_25_20_io_out_sum_exp),
    .io_out_kv(local_pes_25_20_io_out_kv),
    .io_out_stage(local_pes_25_20_io_out_stage)
  );
  PE_1 local_pes_25_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_21_clock),
    .reset(local_pes_25_21_reset),
    .io_in_q(local_pes_25_21_io_in_q),
    .io_in_sum(local_pes_25_21_io_in_sum),
    .io_in_sum_exp(local_pes_25_21_io_in_sum_exp),
    .io_in_kv(local_pes_25_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_21_io_in_inv_sum),
    .io_in_stage(local_pes_25_21_io_in_stage),
    .io_out_q(local_pes_25_21_io_out_q),
    .io_out_sum(local_pes_25_21_io_out_sum),
    .io_out_sum_exp(local_pes_25_21_io_out_sum_exp),
    .io_out_kv(local_pes_25_21_io_out_kv),
    .io_out_stage(local_pes_25_21_io_out_stage)
  );
  PE_1 local_pes_25_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_22_clock),
    .reset(local_pes_25_22_reset),
    .io_in_q(local_pes_25_22_io_in_q),
    .io_in_sum(local_pes_25_22_io_in_sum),
    .io_in_sum_exp(local_pes_25_22_io_in_sum_exp),
    .io_in_kv(local_pes_25_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_22_io_in_inv_sum),
    .io_in_stage(local_pes_25_22_io_in_stage),
    .io_out_q(local_pes_25_22_io_out_q),
    .io_out_sum(local_pes_25_22_io_out_sum),
    .io_out_sum_exp(local_pes_25_22_io_out_sum_exp),
    .io_out_kv(local_pes_25_22_io_out_kv),
    .io_out_stage(local_pes_25_22_io_out_stage)
  );
  PE_1 local_pes_25_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_23_clock),
    .reset(local_pes_25_23_reset),
    .io_in_q(local_pes_25_23_io_in_q),
    .io_in_sum(local_pes_25_23_io_in_sum),
    .io_in_sum_exp(local_pes_25_23_io_in_sum_exp),
    .io_in_kv(local_pes_25_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_23_io_in_inv_sum),
    .io_in_stage(local_pes_25_23_io_in_stage),
    .io_out_q(local_pes_25_23_io_out_q),
    .io_out_sum(local_pes_25_23_io_out_sum),
    .io_out_sum_exp(local_pes_25_23_io_out_sum_exp),
    .io_out_kv(local_pes_25_23_io_out_kv),
    .io_out_stage(local_pes_25_23_io_out_stage)
  );
  PE_1 local_pes_25_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_24_clock),
    .reset(local_pes_25_24_reset),
    .io_in_q(local_pes_25_24_io_in_q),
    .io_in_sum(local_pes_25_24_io_in_sum),
    .io_in_sum_exp(local_pes_25_24_io_in_sum_exp),
    .io_in_kv(local_pes_25_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_24_io_in_inv_sum),
    .io_in_stage(local_pes_25_24_io_in_stage),
    .io_out_q(local_pes_25_24_io_out_q),
    .io_out_sum(local_pes_25_24_io_out_sum),
    .io_out_sum_exp(local_pes_25_24_io_out_sum_exp),
    .io_out_kv(local_pes_25_24_io_out_kv),
    .io_out_stage(local_pes_25_24_io_out_stage)
  );
  PE_1 local_pes_25_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_25_clock),
    .reset(local_pes_25_25_reset),
    .io_in_q(local_pes_25_25_io_in_q),
    .io_in_sum(local_pes_25_25_io_in_sum),
    .io_in_sum_exp(local_pes_25_25_io_in_sum_exp),
    .io_in_kv(local_pes_25_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_25_io_in_inv_sum),
    .io_in_stage(local_pes_25_25_io_in_stage),
    .io_out_q(local_pes_25_25_io_out_q),
    .io_out_sum(local_pes_25_25_io_out_sum),
    .io_out_sum_exp(local_pes_25_25_io_out_sum_exp),
    .io_out_kv(local_pes_25_25_io_out_kv),
    .io_out_stage(local_pes_25_25_io_out_stage)
  );
  PE_1 local_pes_25_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_26_clock),
    .reset(local_pes_25_26_reset),
    .io_in_q(local_pes_25_26_io_in_q),
    .io_in_sum(local_pes_25_26_io_in_sum),
    .io_in_sum_exp(local_pes_25_26_io_in_sum_exp),
    .io_in_kv(local_pes_25_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_26_io_in_inv_sum),
    .io_in_stage(local_pes_25_26_io_in_stage),
    .io_out_q(local_pes_25_26_io_out_q),
    .io_out_sum(local_pes_25_26_io_out_sum),
    .io_out_sum_exp(local_pes_25_26_io_out_sum_exp),
    .io_out_kv(local_pes_25_26_io_out_kv),
    .io_out_stage(local_pes_25_26_io_out_stage)
  );
  PE_1 local_pes_25_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_27_clock),
    .reset(local_pes_25_27_reset),
    .io_in_q(local_pes_25_27_io_in_q),
    .io_in_sum(local_pes_25_27_io_in_sum),
    .io_in_sum_exp(local_pes_25_27_io_in_sum_exp),
    .io_in_kv(local_pes_25_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_27_io_in_inv_sum),
    .io_in_stage(local_pes_25_27_io_in_stage),
    .io_out_q(local_pes_25_27_io_out_q),
    .io_out_sum(local_pes_25_27_io_out_sum),
    .io_out_sum_exp(local_pes_25_27_io_out_sum_exp),
    .io_out_kv(local_pes_25_27_io_out_kv),
    .io_out_stage(local_pes_25_27_io_out_stage)
  );
  PE_1 local_pes_25_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_28_clock),
    .reset(local_pes_25_28_reset),
    .io_in_q(local_pes_25_28_io_in_q),
    .io_in_sum(local_pes_25_28_io_in_sum),
    .io_in_sum_exp(local_pes_25_28_io_in_sum_exp),
    .io_in_kv(local_pes_25_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_28_io_in_inv_sum),
    .io_in_stage(local_pes_25_28_io_in_stage),
    .io_out_q(local_pes_25_28_io_out_q),
    .io_out_sum(local_pes_25_28_io_out_sum),
    .io_out_sum_exp(local_pes_25_28_io_out_sum_exp),
    .io_out_kv(local_pes_25_28_io_out_kv),
    .io_out_stage(local_pes_25_28_io_out_stage)
  );
  PE_1 local_pes_25_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_29_clock),
    .reset(local_pes_25_29_reset),
    .io_in_q(local_pes_25_29_io_in_q),
    .io_in_sum(local_pes_25_29_io_in_sum),
    .io_in_sum_exp(local_pes_25_29_io_in_sum_exp),
    .io_in_kv(local_pes_25_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_29_io_in_inv_sum),
    .io_in_stage(local_pes_25_29_io_in_stage),
    .io_out_q(local_pes_25_29_io_out_q),
    .io_out_sum(local_pes_25_29_io_out_sum),
    .io_out_sum_exp(local_pes_25_29_io_out_sum_exp),
    .io_out_kv(local_pes_25_29_io_out_kv),
    .io_out_stage(local_pes_25_29_io_out_stage)
  );
  PE_1 local_pes_25_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_30_clock),
    .reset(local_pes_25_30_reset),
    .io_in_q(local_pes_25_30_io_in_q),
    .io_in_sum(local_pes_25_30_io_in_sum),
    .io_in_sum_exp(local_pes_25_30_io_in_sum_exp),
    .io_in_kv(local_pes_25_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_30_io_in_inv_sum),
    .io_in_stage(local_pes_25_30_io_in_stage),
    .io_out_q(local_pes_25_30_io_out_q),
    .io_out_sum(local_pes_25_30_io_out_sum),
    .io_out_sum_exp(local_pes_25_30_io_out_sum_exp),
    .io_out_kv(local_pes_25_30_io_out_kv),
    .io_out_stage(local_pes_25_30_io_out_stage)
  );
  PE_1 local_pes_25_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_25_31_clock),
    .reset(local_pes_25_31_reset),
    .io_in_q(local_pes_25_31_io_in_q),
    .io_in_sum(local_pes_25_31_io_in_sum),
    .io_in_sum_exp(local_pes_25_31_io_in_sum_exp),
    .io_in_kv(local_pes_25_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_25_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_25_31_io_in_inv_sum),
    .io_in_stage(local_pes_25_31_io_in_stage),
    .io_out_q(local_pes_25_31_io_out_q),
    .io_out_sum(local_pes_25_31_io_out_sum),
    .io_out_sum_exp(local_pes_25_31_io_out_sum_exp),
    .io_out_kv(local_pes_25_31_io_out_kv),
    .io_out_stage(local_pes_25_31_io_out_stage)
  );
  PE local_pes_26_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_0_clock),
    .reset(local_pes_26_0_reset),
    .io_in_q(local_pes_26_0_io_in_q),
    .io_in_kv(local_pes_26_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_0_io_in_inv_sum),
    .io_in_stage(local_pes_26_0_io_in_stage),
    .io_out_q(local_pes_26_0_io_out_q),
    .io_out_sum(local_pes_26_0_io_out_sum),
    .io_out_kv(local_pes_26_0_io_out_kv),
    .io_out_stage(local_pes_26_0_io_out_stage)
  );
  PE_1 local_pes_26_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_1_clock),
    .reset(local_pes_26_1_reset),
    .io_in_q(local_pes_26_1_io_in_q),
    .io_in_sum(local_pes_26_1_io_in_sum),
    .io_in_sum_exp(local_pes_26_1_io_in_sum_exp),
    .io_in_kv(local_pes_26_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_1_io_in_inv_sum),
    .io_in_stage(local_pes_26_1_io_in_stage),
    .io_out_q(local_pes_26_1_io_out_q),
    .io_out_sum(local_pes_26_1_io_out_sum),
    .io_out_sum_exp(local_pes_26_1_io_out_sum_exp),
    .io_out_kv(local_pes_26_1_io_out_kv),
    .io_out_stage(local_pes_26_1_io_out_stage)
  );
  PE_1 local_pes_26_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_2_clock),
    .reset(local_pes_26_2_reset),
    .io_in_q(local_pes_26_2_io_in_q),
    .io_in_sum(local_pes_26_2_io_in_sum),
    .io_in_sum_exp(local_pes_26_2_io_in_sum_exp),
    .io_in_kv(local_pes_26_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_2_io_in_inv_sum),
    .io_in_stage(local_pes_26_2_io_in_stage),
    .io_out_q(local_pes_26_2_io_out_q),
    .io_out_sum(local_pes_26_2_io_out_sum),
    .io_out_sum_exp(local_pes_26_2_io_out_sum_exp),
    .io_out_kv(local_pes_26_2_io_out_kv),
    .io_out_stage(local_pes_26_2_io_out_stage)
  );
  PE_1 local_pes_26_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_3_clock),
    .reset(local_pes_26_3_reset),
    .io_in_q(local_pes_26_3_io_in_q),
    .io_in_sum(local_pes_26_3_io_in_sum),
    .io_in_sum_exp(local_pes_26_3_io_in_sum_exp),
    .io_in_kv(local_pes_26_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_3_io_in_inv_sum),
    .io_in_stage(local_pes_26_3_io_in_stage),
    .io_out_q(local_pes_26_3_io_out_q),
    .io_out_sum(local_pes_26_3_io_out_sum),
    .io_out_sum_exp(local_pes_26_3_io_out_sum_exp),
    .io_out_kv(local_pes_26_3_io_out_kv),
    .io_out_stage(local_pes_26_3_io_out_stage)
  );
  PE_1 local_pes_26_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_4_clock),
    .reset(local_pes_26_4_reset),
    .io_in_q(local_pes_26_4_io_in_q),
    .io_in_sum(local_pes_26_4_io_in_sum),
    .io_in_sum_exp(local_pes_26_4_io_in_sum_exp),
    .io_in_kv(local_pes_26_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_4_io_in_inv_sum),
    .io_in_stage(local_pes_26_4_io_in_stage),
    .io_out_q(local_pes_26_4_io_out_q),
    .io_out_sum(local_pes_26_4_io_out_sum),
    .io_out_sum_exp(local_pes_26_4_io_out_sum_exp),
    .io_out_kv(local_pes_26_4_io_out_kv),
    .io_out_stage(local_pes_26_4_io_out_stage)
  );
  PE_1 local_pes_26_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_5_clock),
    .reset(local_pes_26_5_reset),
    .io_in_q(local_pes_26_5_io_in_q),
    .io_in_sum(local_pes_26_5_io_in_sum),
    .io_in_sum_exp(local_pes_26_5_io_in_sum_exp),
    .io_in_kv(local_pes_26_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_5_io_in_inv_sum),
    .io_in_stage(local_pes_26_5_io_in_stage),
    .io_out_q(local_pes_26_5_io_out_q),
    .io_out_sum(local_pes_26_5_io_out_sum),
    .io_out_sum_exp(local_pes_26_5_io_out_sum_exp),
    .io_out_kv(local_pes_26_5_io_out_kv),
    .io_out_stage(local_pes_26_5_io_out_stage)
  );
  PE_1 local_pes_26_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_6_clock),
    .reset(local_pes_26_6_reset),
    .io_in_q(local_pes_26_6_io_in_q),
    .io_in_sum(local_pes_26_6_io_in_sum),
    .io_in_sum_exp(local_pes_26_6_io_in_sum_exp),
    .io_in_kv(local_pes_26_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_6_io_in_inv_sum),
    .io_in_stage(local_pes_26_6_io_in_stage),
    .io_out_q(local_pes_26_6_io_out_q),
    .io_out_sum(local_pes_26_6_io_out_sum),
    .io_out_sum_exp(local_pes_26_6_io_out_sum_exp),
    .io_out_kv(local_pes_26_6_io_out_kv),
    .io_out_stage(local_pes_26_6_io_out_stage)
  );
  PE_1 local_pes_26_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_7_clock),
    .reset(local_pes_26_7_reset),
    .io_in_q(local_pes_26_7_io_in_q),
    .io_in_sum(local_pes_26_7_io_in_sum),
    .io_in_sum_exp(local_pes_26_7_io_in_sum_exp),
    .io_in_kv(local_pes_26_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_7_io_in_inv_sum),
    .io_in_stage(local_pes_26_7_io_in_stage),
    .io_out_q(local_pes_26_7_io_out_q),
    .io_out_sum(local_pes_26_7_io_out_sum),
    .io_out_sum_exp(local_pes_26_7_io_out_sum_exp),
    .io_out_kv(local_pes_26_7_io_out_kv),
    .io_out_stage(local_pes_26_7_io_out_stage)
  );
  PE_1 local_pes_26_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_8_clock),
    .reset(local_pes_26_8_reset),
    .io_in_q(local_pes_26_8_io_in_q),
    .io_in_sum(local_pes_26_8_io_in_sum),
    .io_in_sum_exp(local_pes_26_8_io_in_sum_exp),
    .io_in_kv(local_pes_26_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_8_io_in_inv_sum),
    .io_in_stage(local_pes_26_8_io_in_stage),
    .io_out_q(local_pes_26_8_io_out_q),
    .io_out_sum(local_pes_26_8_io_out_sum),
    .io_out_sum_exp(local_pes_26_8_io_out_sum_exp),
    .io_out_kv(local_pes_26_8_io_out_kv),
    .io_out_stage(local_pes_26_8_io_out_stage)
  );
  PE_1 local_pes_26_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_9_clock),
    .reset(local_pes_26_9_reset),
    .io_in_q(local_pes_26_9_io_in_q),
    .io_in_sum(local_pes_26_9_io_in_sum),
    .io_in_sum_exp(local_pes_26_9_io_in_sum_exp),
    .io_in_kv(local_pes_26_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_9_io_in_inv_sum),
    .io_in_stage(local_pes_26_9_io_in_stage),
    .io_out_q(local_pes_26_9_io_out_q),
    .io_out_sum(local_pes_26_9_io_out_sum),
    .io_out_sum_exp(local_pes_26_9_io_out_sum_exp),
    .io_out_kv(local_pes_26_9_io_out_kv),
    .io_out_stage(local_pes_26_9_io_out_stage)
  );
  PE_1 local_pes_26_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_10_clock),
    .reset(local_pes_26_10_reset),
    .io_in_q(local_pes_26_10_io_in_q),
    .io_in_sum(local_pes_26_10_io_in_sum),
    .io_in_sum_exp(local_pes_26_10_io_in_sum_exp),
    .io_in_kv(local_pes_26_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_10_io_in_inv_sum),
    .io_in_stage(local_pes_26_10_io_in_stage),
    .io_out_q(local_pes_26_10_io_out_q),
    .io_out_sum(local_pes_26_10_io_out_sum),
    .io_out_sum_exp(local_pes_26_10_io_out_sum_exp),
    .io_out_kv(local_pes_26_10_io_out_kv),
    .io_out_stage(local_pes_26_10_io_out_stage)
  );
  PE_1 local_pes_26_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_11_clock),
    .reset(local_pes_26_11_reset),
    .io_in_q(local_pes_26_11_io_in_q),
    .io_in_sum(local_pes_26_11_io_in_sum),
    .io_in_sum_exp(local_pes_26_11_io_in_sum_exp),
    .io_in_kv(local_pes_26_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_11_io_in_inv_sum),
    .io_in_stage(local_pes_26_11_io_in_stage),
    .io_out_q(local_pes_26_11_io_out_q),
    .io_out_sum(local_pes_26_11_io_out_sum),
    .io_out_sum_exp(local_pes_26_11_io_out_sum_exp),
    .io_out_kv(local_pes_26_11_io_out_kv),
    .io_out_stage(local_pes_26_11_io_out_stage)
  );
  PE_1 local_pes_26_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_12_clock),
    .reset(local_pes_26_12_reset),
    .io_in_q(local_pes_26_12_io_in_q),
    .io_in_sum(local_pes_26_12_io_in_sum),
    .io_in_sum_exp(local_pes_26_12_io_in_sum_exp),
    .io_in_kv(local_pes_26_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_12_io_in_inv_sum),
    .io_in_stage(local_pes_26_12_io_in_stage),
    .io_out_q(local_pes_26_12_io_out_q),
    .io_out_sum(local_pes_26_12_io_out_sum),
    .io_out_sum_exp(local_pes_26_12_io_out_sum_exp),
    .io_out_kv(local_pes_26_12_io_out_kv),
    .io_out_stage(local_pes_26_12_io_out_stage)
  );
  PE_1 local_pes_26_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_13_clock),
    .reset(local_pes_26_13_reset),
    .io_in_q(local_pes_26_13_io_in_q),
    .io_in_sum(local_pes_26_13_io_in_sum),
    .io_in_sum_exp(local_pes_26_13_io_in_sum_exp),
    .io_in_kv(local_pes_26_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_13_io_in_inv_sum),
    .io_in_stage(local_pes_26_13_io_in_stage),
    .io_out_q(local_pes_26_13_io_out_q),
    .io_out_sum(local_pes_26_13_io_out_sum),
    .io_out_sum_exp(local_pes_26_13_io_out_sum_exp),
    .io_out_kv(local_pes_26_13_io_out_kv),
    .io_out_stage(local_pes_26_13_io_out_stage)
  );
  PE_1 local_pes_26_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_14_clock),
    .reset(local_pes_26_14_reset),
    .io_in_q(local_pes_26_14_io_in_q),
    .io_in_sum(local_pes_26_14_io_in_sum),
    .io_in_sum_exp(local_pes_26_14_io_in_sum_exp),
    .io_in_kv(local_pes_26_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_14_io_in_inv_sum),
    .io_in_stage(local_pes_26_14_io_in_stage),
    .io_out_q(local_pes_26_14_io_out_q),
    .io_out_sum(local_pes_26_14_io_out_sum),
    .io_out_sum_exp(local_pes_26_14_io_out_sum_exp),
    .io_out_kv(local_pes_26_14_io_out_kv),
    .io_out_stage(local_pes_26_14_io_out_stage)
  );
  PE_1 local_pes_26_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_15_clock),
    .reset(local_pes_26_15_reset),
    .io_in_q(local_pes_26_15_io_in_q),
    .io_in_sum(local_pes_26_15_io_in_sum),
    .io_in_sum_exp(local_pes_26_15_io_in_sum_exp),
    .io_in_kv(local_pes_26_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_15_io_in_inv_sum),
    .io_in_stage(local_pes_26_15_io_in_stage),
    .io_out_q(local_pes_26_15_io_out_q),
    .io_out_sum(local_pes_26_15_io_out_sum),
    .io_out_sum_exp(local_pes_26_15_io_out_sum_exp),
    .io_out_kv(local_pes_26_15_io_out_kv),
    .io_out_stage(local_pes_26_15_io_out_stage)
  );
  PE_1 local_pes_26_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_16_clock),
    .reset(local_pes_26_16_reset),
    .io_in_q(local_pes_26_16_io_in_q),
    .io_in_sum(local_pes_26_16_io_in_sum),
    .io_in_sum_exp(local_pes_26_16_io_in_sum_exp),
    .io_in_kv(local_pes_26_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_16_io_in_inv_sum),
    .io_in_stage(local_pes_26_16_io_in_stage),
    .io_out_q(local_pes_26_16_io_out_q),
    .io_out_sum(local_pes_26_16_io_out_sum),
    .io_out_sum_exp(local_pes_26_16_io_out_sum_exp),
    .io_out_kv(local_pes_26_16_io_out_kv),
    .io_out_stage(local_pes_26_16_io_out_stage)
  );
  PE_1 local_pes_26_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_17_clock),
    .reset(local_pes_26_17_reset),
    .io_in_q(local_pes_26_17_io_in_q),
    .io_in_sum(local_pes_26_17_io_in_sum),
    .io_in_sum_exp(local_pes_26_17_io_in_sum_exp),
    .io_in_kv(local_pes_26_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_17_io_in_inv_sum),
    .io_in_stage(local_pes_26_17_io_in_stage),
    .io_out_q(local_pes_26_17_io_out_q),
    .io_out_sum(local_pes_26_17_io_out_sum),
    .io_out_sum_exp(local_pes_26_17_io_out_sum_exp),
    .io_out_kv(local_pes_26_17_io_out_kv),
    .io_out_stage(local_pes_26_17_io_out_stage)
  );
  PE_1 local_pes_26_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_18_clock),
    .reset(local_pes_26_18_reset),
    .io_in_q(local_pes_26_18_io_in_q),
    .io_in_sum(local_pes_26_18_io_in_sum),
    .io_in_sum_exp(local_pes_26_18_io_in_sum_exp),
    .io_in_kv(local_pes_26_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_18_io_in_inv_sum),
    .io_in_stage(local_pes_26_18_io_in_stage),
    .io_out_q(local_pes_26_18_io_out_q),
    .io_out_sum(local_pes_26_18_io_out_sum),
    .io_out_sum_exp(local_pes_26_18_io_out_sum_exp),
    .io_out_kv(local_pes_26_18_io_out_kv),
    .io_out_stage(local_pes_26_18_io_out_stage)
  );
  PE_1 local_pes_26_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_19_clock),
    .reset(local_pes_26_19_reset),
    .io_in_q(local_pes_26_19_io_in_q),
    .io_in_sum(local_pes_26_19_io_in_sum),
    .io_in_sum_exp(local_pes_26_19_io_in_sum_exp),
    .io_in_kv(local_pes_26_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_19_io_in_inv_sum),
    .io_in_stage(local_pes_26_19_io_in_stage),
    .io_out_q(local_pes_26_19_io_out_q),
    .io_out_sum(local_pes_26_19_io_out_sum),
    .io_out_sum_exp(local_pes_26_19_io_out_sum_exp),
    .io_out_kv(local_pes_26_19_io_out_kv),
    .io_out_stage(local_pes_26_19_io_out_stage)
  );
  PE_1 local_pes_26_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_20_clock),
    .reset(local_pes_26_20_reset),
    .io_in_q(local_pes_26_20_io_in_q),
    .io_in_sum(local_pes_26_20_io_in_sum),
    .io_in_sum_exp(local_pes_26_20_io_in_sum_exp),
    .io_in_kv(local_pes_26_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_20_io_in_inv_sum),
    .io_in_stage(local_pes_26_20_io_in_stage),
    .io_out_q(local_pes_26_20_io_out_q),
    .io_out_sum(local_pes_26_20_io_out_sum),
    .io_out_sum_exp(local_pes_26_20_io_out_sum_exp),
    .io_out_kv(local_pes_26_20_io_out_kv),
    .io_out_stage(local_pes_26_20_io_out_stage)
  );
  PE_1 local_pes_26_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_21_clock),
    .reset(local_pes_26_21_reset),
    .io_in_q(local_pes_26_21_io_in_q),
    .io_in_sum(local_pes_26_21_io_in_sum),
    .io_in_sum_exp(local_pes_26_21_io_in_sum_exp),
    .io_in_kv(local_pes_26_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_21_io_in_inv_sum),
    .io_in_stage(local_pes_26_21_io_in_stage),
    .io_out_q(local_pes_26_21_io_out_q),
    .io_out_sum(local_pes_26_21_io_out_sum),
    .io_out_sum_exp(local_pes_26_21_io_out_sum_exp),
    .io_out_kv(local_pes_26_21_io_out_kv),
    .io_out_stage(local_pes_26_21_io_out_stage)
  );
  PE_1 local_pes_26_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_22_clock),
    .reset(local_pes_26_22_reset),
    .io_in_q(local_pes_26_22_io_in_q),
    .io_in_sum(local_pes_26_22_io_in_sum),
    .io_in_sum_exp(local_pes_26_22_io_in_sum_exp),
    .io_in_kv(local_pes_26_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_22_io_in_inv_sum),
    .io_in_stage(local_pes_26_22_io_in_stage),
    .io_out_q(local_pes_26_22_io_out_q),
    .io_out_sum(local_pes_26_22_io_out_sum),
    .io_out_sum_exp(local_pes_26_22_io_out_sum_exp),
    .io_out_kv(local_pes_26_22_io_out_kv),
    .io_out_stage(local_pes_26_22_io_out_stage)
  );
  PE_1 local_pes_26_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_23_clock),
    .reset(local_pes_26_23_reset),
    .io_in_q(local_pes_26_23_io_in_q),
    .io_in_sum(local_pes_26_23_io_in_sum),
    .io_in_sum_exp(local_pes_26_23_io_in_sum_exp),
    .io_in_kv(local_pes_26_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_23_io_in_inv_sum),
    .io_in_stage(local_pes_26_23_io_in_stage),
    .io_out_q(local_pes_26_23_io_out_q),
    .io_out_sum(local_pes_26_23_io_out_sum),
    .io_out_sum_exp(local_pes_26_23_io_out_sum_exp),
    .io_out_kv(local_pes_26_23_io_out_kv),
    .io_out_stage(local_pes_26_23_io_out_stage)
  );
  PE_1 local_pes_26_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_24_clock),
    .reset(local_pes_26_24_reset),
    .io_in_q(local_pes_26_24_io_in_q),
    .io_in_sum(local_pes_26_24_io_in_sum),
    .io_in_sum_exp(local_pes_26_24_io_in_sum_exp),
    .io_in_kv(local_pes_26_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_24_io_in_inv_sum),
    .io_in_stage(local_pes_26_24_io_in_stage),
    .io_out_q(local_pes_26_24_io_out_q),
    .io_out_sum(local_pes_26_24_io_out_sum),
    .io_out_sum_exp(local_pes_26_24_io_out_sum_exp),
    .io_out_kv(local_pes_26_24_io_out_kv),
    .io_out_stage(local_pes_26_24_io_out_stage)
  );
  PE_1 local_pes_26_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_25_clock),
    .reset(local_pes_26_25_reset),
    .io_in_q(local_pes_26_25_io_in_q),
    .io_in_sum(local_pes_26_25_io_in_sum),
    .io_in_sum_exp(local_pes_26_25_io_in_sum_exp),
    .io_in_kv(local_pes_26_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_25_io_in_inv_sum),
    .io_in_stage(local_pes_26_25_io_in_stage),
    .io_out_q(local_pes_26_25_io_out_q),
    .io_out_sum(local_pes_26_25_io_out_sum),
    .io_out_sum_exp(local_pes_26_25_io_out_sum_exp),
    .io_out_kv(local_pes_26_25_io_out_kv),
    .io_out_stage(local_pes_26_25_io_out_stage)
  );
  PE_1 local_pes_26_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_26_clock),
    .reset(local_pes_26_26_reset),
    .io_in_q(local_pes_26_26_io_in_q),
    .io_in_sum(local_pes_26_26_io_in_sum),
    .io_in_sum_exp(local_pes_26_26_io_in_sum_exp),
    .io_in_kv(local_pes_26_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_26_io_in_inv_sum),
    .io_in_stage(local_pes_26_26_io_in_stage),
    .io_out_q(local_pes_26_26_io_out_q),
    .io_out_sum(local_pes_26_26_io_out_sum),
    .io_out_sum_exp(local_pes_26_26_io_out_sum_exp),
    .io_out_kv(local_pes_26_26_io_out_kv),
    .io_out_stage(local_pes_26_26_io_out_stage)
  );
  PE_1 local_pes_26_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_27_clock),
    .reset(local_pes_26_27_reset),
    .io_in_q(local_pes_26_27_io_in_q),
    .io_in_sum(local_pes_26_27_io_in_sum),
    .io_in_sum_exp(local_pes_26_27_io_in_sum_exp),
    .io_in_kv(local_pes_26_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_27_io_in_inv_sum),
    .io_in_stage(local_pes_26_27_io_in_stage),
    .io_out_q(local_pes_26_27_io_out_q),
    .io_out_sum(local_pes_26_27_io_out_sum),
    .io_out_sum_exp(local_pes_26_27_io_out_sum_exp),
    .io_out_kv(local_pes_26_27_io_out_kv),
    .io_out_stage(local_pes_26_27_io_out_stage)
  );
  PE_1 local_pes_26_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_28_clock),
    .reset(local_pes_26_28_reset),
    .io_in_q(local_pes_26_28_io_in_q),
    .io_in_sum(local_pes_26_28_io_in_sum),
    .io_in_sum_exp(local_pes_26_28_io_in_sum_exp),
    .io_in_kv(local_pes_26_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_28_io_in_inv_sum),
    .io_in_stage(local_pes_26_28_io_in_stage),
    .io_out_q(local_pes_26_28_io_out_q),
    .io_out_sum(local_pes_26_28_io_out_sum),
    .io_out_sum_exp(local_pes_26_28_io_out_sum_exp),
    .io_out_kv(local_pes_26_28_io_out_kv),
    .io_out_stage(local_pes_26_28_io_out_stage)
  );
  PE_1 local_pes_26_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_29_clock),
    .reset(local_pes_26_29_reset),
    .io_in_q(local_pes_26_29_io_in_q),
    .io_in_sum(local_pes_26_29_io_in_sum),
    .io_in_sum_exp(local_pes_26_29_io_in_sum_exp),
    .io_in_kv(local_pes_26_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_29_io_in_inv_sum),
    .io_in_stage(local_pes_26_29_io_in_stage),
    .io_out_q(local_pes_26_29_io_out_q),
    .io_out_sum(local_pes_26_29_io_out_sum),
    .io_out_sum_exp(local_pes_26_29_io_out_sum_exp),
    .io_out_kv(local_pes_26_29_io_out_kv),
    .io_out_stage(local_pes_26_29_io_out_stage)
  );
  PE_1 local_pes_26_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_30_clock),
    .reset(local_pes_26_30_reset),
    .io_in_q(local_pes_26_30_io_in_q),
    .io_in_sum(local_pes_26_30_io_in_sum),
    .io_in_sum_exp(local_pes_26_30_io_in_sum_exp),
    .io_in_kv(local_pes_26_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_30_io_in_inv_sum),
    .io_in_stage(local_pes_26_30_io_in_stage),
    .io_out_q(local_pes_26_30_io_out_q),
    .io_out_sum(local_pes_26_30_io_out_sum),
    .io_out_sum_exp(local_pes_26_30_io_out_sum_exp),
    .io_out_kv(local_pes_26_30_io_out_kv),
    .io_out_stage(local_pes_26_30_io_out_stage)
  );
  PE_1 local_pes_26_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_26_31_clock),
    .reset(local_pes_26_31_reset),
    .io_in_q(local_pes_26_31_io_in_q),
    .io_in_sum(local_pes_26_31_io_in_sum),
    .io_in_sum_exp(local_pes_26_31_io_in_sum_exp),
    .io_in_kv(local_pes_26_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_26_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_26_31_io_in_inv_sum),
    .io_in_stage(local_pes_26_31_io_in_stage),
    .io_out_q(local_pes_26_31_io_out_q),
    .io_out_sum(local_pes_26_31_io_out_sum),
    .io_out_sum_exp(local_pes_26_31_io_out_sum_exp),
    .io_out_kv(local_pes_26_31_io_out_kv),
    .io_out_stage(local_pes_26_31_io_out_stage)
  );
  PE local_pes_27_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_0_clock),
    .reset(local_pes_27_0_reset),
    .io_in_q(local_pes_27_0_io_in_q),
    .io_in_kv(local_pes_27_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_0_io_in_inv_sum),
    .io_in_stage(local_pes_27_0_io_in_stage),
    .io_out_q(local_pes_27_0_io_out_q),
    .io_out_sum(local_pes_27_0_io_out_sum),
    .io_out_kv(local_pes_27_0_io_out_kv),
    .io_out_stage(local_pes_27_0_io_out_stage)
  );
  PE_1 local_pes_27_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_1_clock),
    .reset(local_pes_27_1_reset),
    .io_in_q(local_pes_27_1_io_in_q),
    .io_in_sum(local_pes_27_1_io_in_sum),
    .io_in_sum_exp(local_pes_27_1_io_in_sum_exp),
    .io_in_kv(local_pes_27_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_1_io_in_inv_sum),
    .io_in_stage(local_pes_27_1_io_in_stage),
    .io_out_q(local_pes_27_1_io_out_q),
    .io_out_sum(local_pes_27_1_io_out_sum),
    .io_out_sum_exp(local_pes_27_1_io_out_sum_exp),
    .io_out_kv(local_pes_27_1_io_out_kv),
    .io_out_stage(local_pes_27_1_io_out_stage)
  );
  PE_1 local_pes_27_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_2_clock),
    .reset(local_pes_27_2_reset),
    .io_in_q(local_pes_27_2_io_in_q),
    .io_in_sum(local_pes_27_2_io_in_sum),
    .io_in_sum_exp(local_pes_27_2_io_in_sum_exp),
    .io_in_kv(local_pes_27_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_2_io_in_inv_sum),
    .io_in_stage(local_pes_27_2_io_in_stage),
    .io_out_q(local_pes_27_2_io_out_q),
    .io_out_sum(local_pes_27_2_io_out_sum),
    .io_out_sum_exp(local_pes_27_2_io_out_sum_exp),
    .io_out_kv(local_pes_27_2_io_out_kv),
    .io_out_stage(local_pes_27_2_io_out_stage)
  );
  PE_1 local_pes_27_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_3_clock),
    .reset(local_pes_27_3_reset),
    .io_in_q(local_pes_27_3_io_in_q),
    .io_in_sum(local_pes_27_3_io_in_sum),
    .io_in_sum_exp(local_pes_27_3_io_in_sum_exp),
    .io_in_kv(local_pes_27_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_3_io_in_inv_sum),
    .io_in_stage(local_pes_27_3_io_in_stage),
    .io_out_q(local_pes_27_3_io_out_q),
    .io_out_sum(local_pes_27_3_io_out_sum),
    .io_out_sum_exp(local_pes_27_3_io_out_sum_exp),
    .io_out_kv(local_pes_27_3_io_out_kv),
    .io_out_stage(local_pes_27_3_io_out_stage)
  );
  PE_1 local_pes_27_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_4_clock),
    .reset(local_pes_27_4_reset),
    .io_in_q(local_pes_27_4_io_in_q),
    .io_in_sum(local_pes_27_4_io_in_sum),
    .io_in_sum_exp(local_pes_27_4_io_in_sum_exp),
    .io_in_kv(local_pes_27_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_4_io_in_inv_sum),
    .io_in_stage(local_pes_27_4_io_in_stage),
    .io_out_q(local_pes_27_4_io_out_q),
    .io_out_sum(local_pes_27_4_io_out_sum),
    .io_out_sum_exp(local_pes_27_4_io_out_sum_exp),
    .io_out_kv(local_pes_27_4_io_out_kv),
    .io_out_stage(local_pes_27_4_io_out_stage)
  );
  PE_1 local_pes_27_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_5_clock),
    .reset(local_pes_27_5_reset),
    .io_in_q(local_pes_27_5_io_in_q),
    .io_in_sum(local_pes_27_5_io_in_sum),
    .io_in_sum_exp(local_pes_27_5_io_in_sum_exp),
    .io_in_kv(local_pes_27_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_5_io_in_inv_sum),
    .io_in_stage(local_pes_27_5_io_in_stage),
    .io_out_q(local_pes_27_5_io_out_q),
    .io_out_sum(local_pes_27_5_io_out_sum),
    .io_out_sum_exp(local_pes_27_5_io_out_sum_exp),
    .io_out_kv(local_pes_27_5_io_out_kv),
    .io_out_stage(local_pes_27_5_io_out_stage)
  );
  PE_1 local_pes_27_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_6_clock),
    .reset(local_pes_27_6_reset),
    .io_in_q(local_pes_27_6_io_in_q),
    .io_in_sum(local_pes_27_6_io_in_sum),
    .io_in_sum_exp(local_pes_27_6_io_in_sum_exp),
    .io_in_kv(local_pes_27_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_6_io_in_inv_sum),
    .io_in_stage(local_pes_27_6_io_in_stage),
    .io_out_q(local_pes_27_6_io_out_q),
    .io_out_sum(local_pes_27_6_io_out_sum),
    .io_out_sum_exp(local_pes_27_6_io_out_sum_exp),
    .io_out_kv(local_pes_27_6_io_out_kv),
    .io_out_stage(local_pes_27_6_io_out_stage)
  );
  PE_1 local_pes_27_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_7_clock),
    .reset(local_pes_27_7_reset),
    .io_in_q(local_pes_27_7_io_in_q),
    .io_in_sum(local_pes_27_7_io_in_sum),
    .io_in_sum_exp(local_pes_27_7_io_in_sum_exp),
    .io_in_kv(local_pes_27_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_7_io_in_inv_sum),
    .io_in_stage(local_pes_27_7_io_in_stage),
    .io_out_q(local_pes_27_7_io_out_q),
    .io_out_sum(local_pes_27_7_io_out_sum),
    .io_out_sum_exp(local_pes_27_7_io_out_sum_exp),
    .io_out_kv(local_pes_27_7_io_out_kv),
    .io_out_stage(local_pes_27_7_io_out_stage)
  );
  PE_1 local_pes_27_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_8_clock),
    .reset(local_pes_27_8_reset),
    .io_in_q(local_pes_27_8_io_in_q),
    .io_in_sum(local_pes_27_8_io_in_sum),
    .io_in_sum_exp(local_pes_27_8_io_in_sum_exp),
    .io_in_kv(local_pes_27_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_8_io_in_inv_sum),
    .io_in_stage(local_pes_27_8_io_in_stage),
    .io_out_q(local_pes_27_8_io_out_q),
    .io_out_sum(local_pes_27_8_io_out_sum),
    .io_out_sum_exp(local_pes_27_8_io_out_sum_exp),
    .io_out_kv(local_pes_27_8_io_out_kv),
    .io_out_stage(local_pes_27_8_io_out_stage)
  );
  PE_1 local_pes_27_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_9_clock),
    .reset(local_pes_27_9_reset),
    .io_in_q(local_pes_27_9_io_in_q),
    .io_in_sum(local_pes_27_9_io_in_sum),
    .io_in_sum_exp(local_pes_27_9_io_in_sum_exp),
    .io_in_kv(local_pes_27_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_9_io_in_inv_sum),
    .io_in_stage(local_pes_27_9_io_in_stage),
    .io_out_q(local_pes_27_9_io_out_q),
    .io_out_sum(local_pes_27_9_io_out_sum),
    .io_out_sum_exp(local_pes_27_9_io_out_sum_exp),
    .io_out_kv(local_pes_27_9_io_out_kv),
    .io_out_stage(local_pes_27_9_io_out_stage)
  );
  PE_1 local_pes_27_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_10_clock),
    .reset(local_pes_27_10_reset),
    .io_in_q(local_pes_27_10_io_in_q),
    .io_in_sum(local_pes_27_10_io_in_sum),
    .io_in_sum_exp(local_pes_27_10_io_in_sum_exp),
    .io_in_kv(local_pes_27_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_10_io_in_inv_sum),
    .io_in_stage(local_pes_27_10_io_in_stage),
    .io_out_q(local_pes_27_10_io_out_q),
    .io_out_sum(local_pes_27_10_io_out_sum),
    .io_out_sum_exp(local_pes_27_10_io_out_sum_exp),
    .io_out_kv(local_pes_27_10_io_out_kv),
    .io_out_stage(local_pes_27_10_io_out_stage)
  );
  PE_1 local_pes_27_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_11_clock),
    .reset(local_pes_27_11_reset),
    .io_in_q(local_pes_27_11_io_in_q),
    .io_in_sum(local_pes_27_11_io_in_sum),
    .io_in_sum_exp(local_pes_27_11_io_in_sum_exp),
    .io_in_kv(local_pes_27_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_11_io_in_inv_sum),
    .io_in_stage(local_pes_27_11_io_in_stage),
    .io_out_q(local_pes_27_11_io_out_q),
    .io_out_sum(local_pes_27_11_io_out_sum),
    .io_out_sum_exp(local_pes_27_11_io_out_sum_exp),
    .io_out_kv(local_pes_27_11_io_out_kv),
    .io_out_stage(local_pes_27_11_io_out_stage)
  );
  PE_1 local_pes_27_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_12_clock),
    .reset(local_pes_27_12_reset),
    .io_in_q(local_pes_27_12_io_in_q),
    .io_in_sum(local_pes_27_12_io_in_sum),
    .io_in_sum_exp(local_pes_27_12_io_in_sum_exp),
    .io_in_kv(local_pes_27_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_12_io_in_inv_sum),
    .io_in_stage(local_pes_27_12_io_in_stage),
    .io_out_q(local_pes_27_12_io_out_q),
    .io_out_sum(local_pes_27_12_io_out_sum),
    .io_out_sum_exp(local_pes_27_12_io_out_sum_exp),
    .io_out_kv(local_pes_27_12_io_out_kv),
    .io_out_stage(local_pes_27_12_io_out_stage)
  );
  PE_1 local_pes_27_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_13_clock),
    .reset(local_pes_27_13_reset),
    .io_in_q(local_pes_27_13_io_in_q),
    .io_in_sum(local_pes_27_13_io_in_sum),
    .io_in_sum_exp(local_pes_27_13_io_in_sum_exp),
    .io_in_kv(local_pes_27_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_13_io_in_inv_sum),
    .io_in_stage(local_pes_27_13_io_in_stage),
    .io_out_q(local_pes_27_13_io_out_q),
    .io_out_sum(local_pes_27_13_io_out_sum),
    .io_out_sum_exp(local_pes_27_13_io_out_sum_exp),
    .io_out_kv(local_pes_27_13_io_out_kv),
    .io_out_stage(local_pes_27_13_io_out_stage)
  );
  PE_1 local_pes_27_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_14_clock),
    .reset(local_pes_27_14_reset),
    .io_in_q(local_pes_27_14_io_in_q),
    .io_in_sum(local_pes_27_14_io_in_sum),
    .io_in_sum_exp(local_pes_27_14_io_in_sum_exp),
    .io_in_kv(local_pes_27_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_14_io_in_inv_sum),
    .io_in_stage(local_pes_27_14_io_in_stage),
    .io_out_q(local_pes_27_14_io_out_q),
    .io_out_sum(local_pes_27_14_io_out_sum),
    .io_out_sum_exp(local_pes_27_14_io_out_sum_exp),
    .io_out_kv(local_pes_27_14_io_out_kv),
    .io_out_stage(local_pes_27_14_io_out_stage)
  );
  PE_1 local_pes_27_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_15_clock),
    .reset(local_pes_27_15_reset),
    .io_in_q(local_pes_27_15_io_in_q),
    .io_in_sum(local_pes_27_15_io_in_sum),
    .io_in_sum_exp(local_pes_27_15_io_in_sum_exp),
    .io_in_kv(local_pes_27_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_15_io_in_inv_sum),
    .io_in_stage(local_pes_27_15_io_in_stage),
    .io_out_q(local_pes_27_15_io_out_q),
    .io_out_sum(local_pes_27_15_io_out_sum),
    .io_out_sum_exp(local_pes_27_15_io_out_sum_exp),
    .io_out_kv(local_pes_27_15_io_out_kv),
    .io_out_stage(local_pes_27_15_io_out_stage)
  );
  PE_1 local_pes_27_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_16_clock),
    .reset(local_pes_27_16_reset),
    .io_in_q(local_pes_27_16_io_in_q),
    .io_in_sum(local_pes_27_16_io_in_sum),
    .io_in_sum_exp(local_pes_27_16_io_in_sum_exp),
    .io_in_kv(local_pes_27_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_16_io_in_inv_sum),
    .io_in_stage(local_pes_27_16_io_in_stage),
    .io_out_q(local_pes_27_16_io_out_q),
    .io_out_sum(local_pes_27_16_io_out_sum),
    .io_out_sum_exp(local_pes_27_16_io_out_sum_exp),
    .io_out_kv(local_pes_27_16_io_out_kv),
    .io_out_stage(local_pes_27_16_io_out_stage)
  );
  PE_1 local_pes_27_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_17_clock),
    .reset(local_pes_27_17_reset),
    .io_in_q(local_pes_27_17_io_in_q),
    .io_in_sum(local_pes_27_17_io_in_sum),
    .io_in_sum_exp(local_pes_27_17_io_in_sum_exp),
    .io_in_kv(local_pes_27_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_17_io_in_inv_sum),
    .io_in_stage(local_pes_27_17_io_in_stage),
    .io_out_q(local_pes_27_17_io_out_q),
    .io_out_sum(local_pes_27_17_io_out_sum),
    .io_out_sum_exp(local_pes_27_17_io_out_sum_exp),
    .io_out_kv(local_pes_27_17_io_out_kv),
    .io_out_stage(local_pes_27_17_io_out_stage)
  );
  PE_1 local_pes_27_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_18_clock),
    .reset(local_pes_27_18_reset),
    .io_in_q(local_pes_27_18_io_in_q),
    .io_in_sum(local_pes_27_18_io_in_sum),
    .io_in_sum_exp(local_pes_27_18_io_in_sum_exp),
    .io_in_kv(local_pes_27_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_18_io_in_inv_sum),
    .io_in_stage(local_pes_27_18_io_in_stage),
    .io_out_q(local_pes_27_18_io_out_q),
    .io_out_sum(local_pes_27_18_io_out_sum),
    .io_out_sum_exp(local_pes_27_18_io_out_sum_exp),
    .io_out_kv(local_pes_27_18_io_out_kv),
    .io_out_stage(local_pes_27_18_io_out_stage)
  );
  PE_1 local_pes_27_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_19_clock),
    .reset(local_pes_27_19_reset),
    .io_in_q(local_pes_27_19_io_in_q),
    .io_in_sum(local_pes_27_19_io_in_sum),
    .io_in_sum_exp(local_pes_27_19_io_in_sum_exp),
    .io_in_kv(local_pes_27_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_19_io_in_inv_sum),
    .io_in_stage(local_pes_27_19_io_in_stage),
    .io_out_q(local_pes_27_19_io_out_q),
    .io_out_sum(local_pes_27_19_io_out_sum),
    .io_out_sum_exp(local_pes_27_19_io_out_sum_exp),
    .io_out_kv(local_pes_27_19_io_out_kv),
    .io_out_stage(local_pes_27_19_io_out_stage)
  );
  PE_1 local_pes_27_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_20_clock),
    .reset(local_pes_27_20_reset),
    .io_in_q(local_pes_27_20_io_in_q),
    .io_in_sum(local_pes_27_20_io_in_sum),
    .io_in_sum_exp(local_pes_27_20_io_in_sum_exp),
    .io_in_kv(local_pes_27_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_20_io_in_inv_sum),
    .io_in_stage(local_pes_27_20_io_in_stage),
    .io_out_q(local_pes_27_20_io_out_q),
    .io_out_sum(local_pes_27_20_io_out_sum),
    .io_out_sum_exp(local_pes_27_20_io_out_sum_exp),
    .io_out_kv(local_pes_27_20_io_out_kv),
    .io_out_stage(local_pes_27_20_io_out_stage)
  );
  PE_1 local_pes_27_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_21_clock),
    .reset(local_pes_27_21_reset),
    .io_in_q(local_pes_27_21_io_in_q),
    .io_in_sum(local_pes_27_21_io_in_sum),
    .io_in_sum_exp(local_pes_27_21_io_in_sum_exp),
    .io_in_kv(local_pes_27_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_21_io_in_inv_sum),
    .io_in_stage(local_pes_27_21_io_in_stage),
    .io_out_q(local_pes_27_21_io_out_q),
    .io_out_sum(local_pes_27_21_io_out_sum),
    .io_out_sum_exp(local_pes_27_21_io_out_sum_exp),
    .io_out_kv(local_pes_27_21_io_out_kv),
    .io_out_stage(local_pes_27_21_io_out_stage)
  );
  PE_1 local_pes_27_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_22_clock),
    .reset(local_pes_27_22_reset),
    .io_in_q(local_pes_27_22_io_in_q),
    .io_in_sum(local_pes_27_22_io_in_sum),
    .io_in_sum_exp(local_pes_27_22_io_in_sum_exp),
    .io_in_kv(local_pes_27_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_22_io_in_inv_sum),
    .io_in_stage(local_pes_27_22_io_in_stage),
    .io_out_q(local_pes_27_22_io_out_q),
    .io_out_sum(local_pes_27_22_io_out_sum),
    .io_out_sum_exp(local_pes_27_22_io_out_sum_exp),
    .io_out_kv(local_pes_27_22_io_out_kv),
    .io_out_stage(local_pes_27_22_io_out_stage)
  );
  PE_1 local_pes_27_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_23_clock),
    .reset(local_pes_27_23_reset),
    .io_in_q(local_pes_27_23_io_in_q),
    .io_in_sum(local_pes_27_23_io_in_sum),
    .io_in_sum_exp(local_pes_27_23_io_in_sum_exp),
    .io_in_kv(local_pes_27_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_23_io_in_inv_sum),
    .io_in_stage(local_pes_27_23_io_in_stage),
    .io_out_q(local_pes_27_23_io_out_q),
    .io_out_sum(local_pes_27_23_io_out_sum),
    .io_out_sum_exp(local_pes_27_23_io_out_sum_exp),
    .io_out_kv(local_pes_27_23_io_out_kv),
    .io_out_stage(local_pes_27_23_io_out_stage)
  );
  PE_1 local_pes_27_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_24_clock),
    .reset(local_pes_27_24_reset),
    .io_in_q(local_pes_27_24_io_in_q),
    .io_in_sum(local_pes_27_24_io_in_sum),
    .io_in_sum_exp(local_pes_27_24_io_in_sum_exp),
    .io_in_kv(local_pes_27_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_24_io_in_inv_sum),
    .io_in_stage(local_pes_27_24_io_in_stage),
    .io_out_q(local_pes_27_24_io_out_q),
    .io_out_sum(local_pes_27_24_io_out_sum),
    .io_out_sum_exp(local_pes_27_24_io_out_sum_exp),
    .io_out_kv(local_pes_27_24_io_out_kv),
    .io_out_stage(local_pes_27_24_io_out_stage)
  );
  PE_1 local_pes_27_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_25_clock),
    .reset(local_pes_27_25_reset),
    .io_in_q(local_pes_27_25_io_in_q),
    .io_in_sum(local_pes_27_25_io_in_sum),
    .io_in_sum_exp(local_pes_27_25_io_in_sum_exp),
    .io_in_kv(local_pes_27_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_25_io_in_inv_sum),
    .io_in_stage(local_pes_27_25_io_in_stage),
    .io_out_q(local_pes_27_25_io_out_q),
    .io_out_sum(local_pes_27_25_io_out_sum),
    .io_out_sum_exp(local_pes_27_25_io_out_sum_exp),
    .io_out_kv(local_pes_27_25_io_out_kv),
    .io_out_stage(local_pes_27_25_io_out_stage)
  );
  PE_1 local_pes_27_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_26_clock),
    .reset(local_pes_27_26_reset),
    .io_in_q(local_pes_27_26_io_in_q),
    .io_in_sum(local_pes_27_26_io_in_sum),
    .io_in_sum_exp(local_pes_27_26_io_in_sum_exp),
    .io_in_kv(local_pes_27_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_26_io_in_inv_sum),
    .io_in_stage(local_pes_27_26_io_in_stage),
    .io_out_q(local_pes_27_26_io_out_q),
    .io_out_sum(local_pes_27_26_io_out_sum),
    .io_out_sum_exp(local_pes_27_26_io_out_sum_exp),
    .io_out_kv(local_pes_27_26_io_out_kv),
    .io_out_stage(local_pes_27_26_io_out_stage)
  );
  PE_1 local_pes_27_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_27_clock),
    .reset(local_pes_27_27_reset),
    .io_in_q(local_pes_27_27_io_in_q),
    .io_in_sum(local_pes_27_27_io_in_sum),
    .io_in_sum_exp(local_pes_27_27_io_in_sum_exp),
    .io_in_kv(local_pes_27_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_27_io_in_inv_sum),
    .io_in_stage(local_pes_27_27_io_in_stage),
    .io_out_q(local_pes_27_27_io_out_q),
    .io_out_sum(local_pes_27_27_io_out_sum),
    .io_out_sum_exp(local_pes_27_27_io_out_sum_exp),
    .io_out_kv(local_pes_27_27_io_out_kv),
    .io_out_stage(local_pes_27_27_io_out_stage)
  );
  PE_1 local_pes_27_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_28_clock),
    .reset(local_pes_27_28_reset),
    .io_in_q(local_pes_27_28_io_in_q),
    .io_in_sum(local_pes_27_28_io_in_sum),
    .io_in_sum_exp(local_pes_27_28_io_in_sum_exp),
    .io_in_kv(local_pes_27_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_28_io_in_inv_sum),
    .io_in_stage(local_pes_27_28_io_in_stage),
    .io_out_q(local_pes_27_28_io_out_q),
    .io_out_sum(local_pes_27_28_io_out_sum),
    .io_out_sum_exp(local_pes_27_28_io_out_sum_exp),
    .io_out_kv(local_pes_27_28_io_out_kv),
    .io_out_stage(local_pes_27_28_io_out_stage)
  );
  PE_1 local_pes_27_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_29_clock),
    .reset(local_pes_27_29_reset),
    .io_in_q(local_pes_27_29_io_in_q),
    .io_in_sum(local_pes_27_29_io_in_sum),
    .io_in_sum_exp(local_pes_27_29_io_in_sum_exp),
    .io_in_kv(local_pes_27_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_29_io_in_inv_sum),
    .io_in_stage(local_pes_27_29_io_in_stage),
    .io_out_q(local_pes_27_29_io_out_q),
    .io_out_sum(local_pes_27_29_io_out_sum),
    .io_out_sum_exp(local_pes_27_29_io_out_sum_exp),
    .io_out_kv(local_pes_27_29_io_out_kv),
    .io_out_stage(local_pes_27_29_io_out_stage)
  );
  PE_1 local_pes_27_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_30_clock),
    .reset(local_pes_27_30_reset),
    .io_in_q(local_pes_27_30_io_in_q),
    .io_in_sum(local_pes_27_30_io_in_sum),
    .io_in_sum_exp(local_pes_27_30_io_in_sum_exp),
    .io_in_kv(local_pes_27_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_30_io_in_inv_sum),
    .io_in_stage(local_pes_27_30_io_in_stage),
    .io_out_q(local_pes_27_30_io_out_q),
    .io_out_sum(local_pes_27_30_io_out_sum),
    .io_out_sum_exp(local_pes_27_30_io_out_sum_exp),
    .io_out_kv(local_pes_27_30_io_out_kv),
    .io_out_stage(local_pes_27_30_io_out_stage)
  );
  PE_1 local_pes_27_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_27_31_clock),
    .reset(local_pes_27_31_reset),
    .io_in_q(local_pes_27_31_io_in_q),
    .io_in_sum(local_pes_27_31_io_in_sum),
    .io_in_sum_exp(local_pes_27_31_io_in_sum_exp),
    .io_in_kv(local_pes_27_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_27_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_27_31_io_in_inv_sum),
    .io_in_stage(local_pes_27_31_io_in_stage),
    .io_out_q(local_pes_27_31_io_out_q),
    .io_out_sum(local_pes_27_31_io_out_sum),
    .io_out_sum_exp(local_pes_27_31_io_out_sum_exp),
    .io_out_kv(local_pes_27_31_io_out_kv),
    .io_out_stage(local_pes_27_31_io_out_stage)
  );
  PE local_pes_28_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_0_clock),
    .reset(local_pes_28_0_reset),
    .io_in_q(local_pes_28_0_io_in_q),
    .io_in_kv(local_pes_28_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_0_io_in_inv_sum),
    .io_in_stage(local_pes_28_0_io_in_stage),
    .io_out_q(local_pes_28_0_io_out_q),
    .io_out_sum(local_pes_28_0_io_out_sum),
    .io_out_kv(local_pes_28_0_io_out_kv),
    .io_out_stage(local_pes_28_0_io_out_stage)
  );
  PE_1 local_pes_28_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_1_clock),
    .reset(local_pes_28_1_reset),
    .io_in_q(local_pes_28_1_io_in_q),
    .io_in_sum(local_pes_28_1_io_in_sum),
    .io_in_sum_exp(local_pes_28_1_io_in_sum_exp),
    .io_in_kv(local_pes_28_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_1_io_in_inv_sum),
    .io_in_stage(local_pes_28_1_io_in_stage),
    .io_out_q(local_pes_28_1_io_out_q),
    .io_out_sum(local_pes_28_1_io_out_sum),
    .io_out_sum_exp(local_pes_28_1_io_out_sum_exp),
    .io_out_kv(local_pes_28_1_io_out_kv),
    .io_out_stage(local_pes_28_1_io_out_stage)
  );
  PE_1 local_pes_28_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_2_clock),
    .reset(local_pes_28_2_reset),
    .io_in_q(local_pes_28_2_io_in_q),
    .io_in_sum(local_pes_28_2_io_in_sum),
    .io_in_sum_exp(local_pes_28_2_io_in_sum_exp),
    .io_in_kv(local_pes_28_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_2_io_in_inv_sum),
    .io_in_stage(local_pes_28_2_io_in_stage),
    .io_out_q(local_pes_28_2_io_out_q),
    .io_out_sum(local_pes_28_2_io_out_sum),
    .io_out_sum_exp(local_pes_28_2_io_out_sum_exp),
    .io_out_kv(local_pes_28_2_io_out_kv),
    .io_out_stage(local_pes_28_2_io_out_stage)
  );
  PE_1 local_pes_28_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_3_clock),
    .reset(local_pes_28_3_reset),
    .io_in_q(local_pes_28_3_io_in_q),
    .io_in_sum(local_pes_28_3_io_in_sum),
    .io_in_sum_exp(local_pes_28_3_io_in_sum_exp),
    .io_in_kv(local_pes_28_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_3_io_in_inv_sum),
    .io_in_stage(local_pes_28_3_io_in_stage),
    .io_out_q(local_pes_28_3_io_out_q),
    .io_out_sum(local_pes_28_3_io_out_sum),
    .io_out_sum_exp(local_pes_28_3_io_out_sum_exp),
    .io_out_kv(local_pes_28_3_io_out_kv),
    .io_out_stage(local_pes_28_3_io_out_stage)
  );
  PE_1 local_pes_28_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_4_clock),
    .reset(local_pes_28_4_reset),
    .io_in_q(local_pes_28_4_io_in_q),
    .io_in_sum(local_pes_28_4_io_in_sum),
    .io_in_sum_exp(local_pes_28_4_io_in_sum_exp),
    .io_in_kv(local_pes_28_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_4_io_in_inv_sum),
    .io_in_stage(local_pes_28_4_io_in_stage),
    .io_out_q(local_pes_28_4_io_out_q),
    .io_out_sum(local_pes_28_4_io_out_sum),
    .io_out_sum_exp(local_pes_28_4_io_out_sum_exp),
    .io_out_kv(local_pes_28_4_io_out_kv),
    .io_out_stage(local_pes_28_4_io_out_stage)
  );
  PE_1 local_pes_28_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_5_clock),
    .reset(local_pes_28_5_reset),
    .io_in_q(local_pes_28_5_io_in_q),
    .io_in_sum(local_pes_28_5_io_in_sum),
    .io_in_sum_exp(local_pes_28_5_io_in_sum_exp),
    .io_in_kv(local_pes_28_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_5_io_in_inv_sum),
    .io_in_stage(local_pes_28_5_io_in_stage),
    .io_out_q(local_pes_28_5_io_out_q),
    .io_out_sum(local_pes_28_5_io_out_sum),
    .io_out_sum_exp(local_pes_28_5_io_out_sum_exp),
    .io_out_kv(local_pes_28_5_io_out_kv),
    .io_out_stage(local_pes_28_5_io_out_stage)
  );
  PE_1 local_pes_28_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_6_clock),
    .reset(local_pes_28_6_reset),
    .io_in_q(local_pes_28_6_io_in_q),
    .io_in_sum(local_pes_28_6_io_in_sum),
    .io_in_sum_exp(local_pes_28_6_io_in_sum_exp),
    .io_in_kv(local_pes_28_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_6_io_in_inv_sum),
    .io_in_stage(local_pes_28_6_io_in_stage),
    .io_out_q(local_pes_28_6_io_out_q),
    .io_out_sum(local_pes_28_6_io_out_sum),
    .io_out_sum_exp(local_pes_28_6_io_out_sum_exp),
    .io_out_kv(local_pes_28_6_io_out_kv),
    .io_out_stage(local_pes_28_6_io_out_stage)
  );
  PE_1 local_pes_28_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_7_clock),
    .reset(local_pes_28_7_reset),
    .io_in_q(local_pes_28_7_io_in_q),
    .io_in_sum(local_pes_28_7_io_in_sum),
    .io_in_sum_exp(local_pes_28_7_io_in_sum_exp),
    .io_in_kv(local_pes_28_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_7_io_in_inv_sum),
    .io_in_stage(local_pes_28_7_io_in_stage),
    .io_out_q(local_pes_28_7_io_out_q),
    .io_out_sum(local_pes_28_7_io_out_sum),
    .io_out_sum_exp(local_pes_28_7_io_out_sum_exp),
    .io_out_kv(local_pes_28_7_io_out_kv),
    .io_out_stage(local_pes_28_7_io_out_stage)
  );
  PE_1 local_pes_28_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_8_clock),
    .reset(local_pes_28_8_reset),
    .io_in_q(local_pes_28_8_io_in_q),
    .io_in_sum(local_pes_28_8_io_in_sum),
    .io_in_sum_exp(local_pes_28_8_io_in_sum_exp),
    .io_in_kv(local_pes_28_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_8_io_in_inv_sum),
    .io_in_stage(local_pes_28_8_io_in_stage),
    .io_out_q(local_pes_28_8_io_out_q),
    .io_out_sum(local_pes_28_8_io_out_sum),
    .io_out_sum_exp(local_pes_28_8_io_out_sum_exp),
    .io_out_kv(local_pes_28_8_io_out_kv),
    .io_out_stage(local_pes_28_8_io_out_stage)
  );
  PE_1 local_pes_28_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_9_clock),
    .reset(local_pes_28_9_reset),
    .io_in_q(local_pes_28_9_io_in_q),
    .io_in_sum(local_pes_28_9_io_in_sum),
    .io_in_sum_exp(local_pes_28_9_io_in_sum_exp),
    .io_in_kv(local_pes_28_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_9_io_in_inv_sum),
    .io_in_stage(local_pes_28_9_io_in_stage),
    .io_out_q(local_pes_28_9_io_out_q),
    .io_out_sum(local_pes_28_9_io_out_sum),
    .io_out_sum_exp(local_pes_28_9_io_out_sum_exp),
    .io_out_kv(local_pes_28_9_io_out_kv),
    .io_out_stage(local_pes_28_9_io_out_stage)
  );
  PE_1 local_pes_28_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_10_clock),
    .reset(local_pes_28_10_reset),
    .io_in_q(local_pes_28_10_io_in_q),
    .io_in_sum(local_pes_28_10_io_in_sum),
    .io_in_sum_exp(local_pes_28_10_io_in_sum_exp),
    .io_in_kv(local_pes_28_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_10_io_in_inv_sum),
    .io_in_stage(local_pes_28_10_io_in_stage),
    .io_out_q(local_pes_28_10_io_out_q),
    .io_out_sum(local_pes_28_10_io_out_sum),
    .io_out_sum_exp(local_pes_28_10_io_out_sum_exp),
    .io_out_kv(local_pes_28_10_io_out_kv),
    .io_out_stage(local_pes_28_10_io_out_stage)
  );
  PE_1 local_pes_28_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_11_clock),
    .reset(local_pes_28_11_reset),
    .io_in_q(local_pes_28_11_io_in_q),
    .io_in_sum(local_pes_28_11_io_in_sum),
    .io_in_sum_exp(local_pes_28_11_io_in_sum_exp),
    .io_in_kv(local_pes_28_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_11_io_in_inv_sum),
    .io_in_stage(local_pes_28_11_io_in_stage),
    .io_out_q(local_pes_28_11_io_out_q),
    .io_out_sum(local_pes_28_11_io_out_sum),
    .io_out_sum_exp(local_pes_28_11_io_out_sum_exp),
    .io_out_kv(local_pes_28_11_io_out_kv),
    .io_out_stage(local_pes_28_11_io_out_stage)
  );
  PE_1 local_pes_28_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_12_clock),
    .reset(local_pes_28_12_reset),
    .io_in_q(local_pes_28_12_io_in_q),
    .io_in_sum(local_pes_28_12_io_in_sum),
    .io_in_sum_exp(local_pes_28_12_io_in_sum_exp),
    .io_in_kv(local_pes_28_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_12_io_in_inv_sum),
    .io_in_stage(local_pes_28_12_io_in_stage),
    .io_out_q(local_pes_28_12_io_out_q),
    .io_out_sum(local_pes_28_12_io_out_sum),
    .io_out_sum_exp(local_pes_28_12_io_out_sum_exp),
    .io_out_kv(local_pes_28_12_io_out_kv),
    .io_out_stage(local_pes_28_12_io_out_stage)
  );
  PE_1 local_pes_28_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_13_clock),
    .reset(local_pes_28_13_reset),
    .io_in_q(local_pes_28_13_io_in_q),
    .io_in_sum(local_pes_28_13_io_in_sum),
    .io_in_sum_exp(local_pes_28_13_io_in_sum_exp),
    .io_in_kv(local_pes_28_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_13_io_in_inv_sum),
    .io_in_stage(local_pes_28_13_io_in_stage),
    .io_out_q(local_pes_28_13_io_out_q),
    .io_out_sum(local_pes_28_13_io_out_sum),
    .io_out_sum_exp(local_pes_28_13_io_out_sum_exp),
    .io_out_kv(local_pes_28_13_io_out_kv),
    .io_out_stage(local_pes_28_13_io_out_stage)
  );
  PE_1 local_pes_28_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_14_clock),
    .reset(local_pes_28_14_reset),
    .io_in_q(local_pes_28_14_io_in_q),
    .io_in_sum(local_pes_28_14_io_in_sum),
    .io_in_sum_exp(local_pes_28_14_io_in_sum_exp),
    .io_in_kv(local_pes_28_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_14_io_in_inv_sum),
    .io_in_stage(local_pes_28_14_io_in_stage),
    .io_out_q(local_pes_28_14_io_out_q),
    .io_out_sum(local_pes_28_14_io_out_sum),
    .io_out_sum_exp(local_pes_28_14_io_out_sum_exp),
    .io_out_kv(local_pes_28_14_io_out_kv),
    .io_out_stage(local_pes_28_14_io_out_stage)
  );
  PE_1 local_pes_28_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_15_clock),
    .reset(local_pes_28_15_reset),
    .io_in_q(local_pes_28_15_io_in_q),
    .io_in_sum(local_pes_28_15_io_in_sum),
    .io_in_sum_exp(local_pes_28_15_io_in_sum_exp),
    .io_in_kv(local_pes_28_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_15_io_in_inv_sum),
    .io_in_stage(local_pes_28_15_io_in_stage),
    .io_out_q(local_pes_28_15_io_out_q),
    .io_out_sum(local_pes_28_15_io_out_sum),
    .io_out_sum_exp(local_pes_28_15_io_out_sum_exp),
    .io_out_kv(local_pes_28_15_io_out_kv),
    .io_out_stage(local_pes_28_15_io_out_stage)
  );
  PE_1 local_pes_28_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_16_clock),
    .reset(local_pes_28_16_reset),
    .io_in_q(local_pes_28_16_io_in_q),
    .io_in_sum(local_pes_28_16_io_in_sum),
    .io_in_sum_exp(local_pes_28_16_io_in_sum_exp),
    .io_in_kv(local_pes_28_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_16_io_in_inv_sum),
    .io_in_stage(local_pes_28_16_io_in_stage),
    .io_out_q(local_pes_28_16_io_out_q),
    .io_out_sum(local_pes_28_16_io_out_sum),
    .io_out_sum_exp(local_pes_28_16_io_out_sum_exp),
    .io_out_kv(local_pes_28_16_io_out_kv),
    .io_out_stage(local_pes_28_16_io_out_stage)
  );
  PE_1 local_pes_28_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_17_clock),
    .reset(local_pes_28_17_reset),
    .io_in_q(local_pes_28_17_io_in_q),
    .io_in_sum(local_pes_28_17_io_in_sum),
    .io_in_sum_exp(local_pes_28_17_io_in_sum_exp),
    .io_in_kv(local_pes_28_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_17_io_in_inv_sum),
    .io_in_stage(local_pes_28_17_io_in_stage),
    .io_out_q(local_pes_28_17_io_out_q),
    .io_out_sum(local_pes_28_17_io_out_sum),
    .io_out_sum_exp(local_pes_28_17_io_out_sum_exp),
    .io_out_kv(local_pes_28_17_io_out_kv),
    .io_out_stage(local_pes_28_17_io_out_stage)
  );
  PE_1 local_pes_28_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_18_clock),
    .reset(local_pes_28_18_reset),
    .io_in_q(local_pes_28_18_io_in_q),
    .io_in_sum(local_pes_28_18_io_in_sum),
    .io_in_sum_exp(local_pes_28_18_io_in_sum_exp),
    .io_in_kv(local_pes_28_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_18_io_in_inv_sum),
    .io_in_stage(local_pes_28_18_io_in_stage),
    .io_out_q(local_pes_28_18_io_out_q),
    .io_out_sum(local_pes_28_18_io_out_sum),
    .io_out_sum_exp(local_pes_28_18_io_out_sum_exp),
    .io_out_kv(local_pes_28_18_io_out_kv),
    .io_out_stage(local_pes_28_18_io_out_stage)
  );
  PE_1 local_pes_28_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_19_clock),
    .reset(local_pes_28_19_reset),
    .io_in_q(local_pes_28_19_io_in_q),
    .io_in_sum(local_pes_28_19_io_in_sum),
    .io_in_sum_exp(local_pes_28_19_io_in_sum_exp),
    .io_in_kv(local_pes_28_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_19_io_in_inv_sum),
    .io_in_stage(local_pes_28_19_io_in_stage),
    .io_out_q(local_pes_28_19_io_out_q),
    .io_out_sum(local_pes_28_19_io_out_sum),
    .io_out_sum_exp(local_pes_28_19_io_out_sum_exp),
    .io_out_kv(local_pes_28_19_io_out_kv),
    .io_out_stage(local_pes_28_19_io_out_stage)
  );
  PE_1 local_pes_28_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_20_clock),
    .reset(local_pes_28_20_reset),
    .io_in_q(local_pes_28_20_io_in_q),
    .io_in_sum(local_pes_28_20_io_in_sum),
    .io_in_sum_exp(local_pes_28_20_io_in_sum_exp),
    .io_in_kv(local_pes_28_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_20_io_in_inv_sum),
    .io_in_stage(local_pes_28_20_io_in_stage),
    .io_out_q(local_pes_28_20_io_out_q),
    .io_out_sum(local_pes_28_20_io_out_sum),
    .io_out_sum_exp(local_pes_28_20_io_out_sum_exp),
    .io_out_kv(local_pes_28_20_io_out_kv),
    .io_out_stage(local_pes_28_20_io_out_stage)
  );
  PE_1 local_pes_28_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_21_clock),
    .reset(local_pes_28_21_reset),
    .io_in_q(local_pes_28_21_io_in_q),
    .io_in_sum(local_pes_28_21_io_in_sum),
    .io_in_sum_exp(local_pes_28_21_io_in_sum_exp),
    .io_in_kv(local_pes_28_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_21_io_in_inv_sum),
    .io_in_stage(local_pes_28_21_io_in_stage),
    .io_out_q(local_pes_28_21_io_out_q),
    .io_out_sum(local_pes_28_21_io_out_sum),
    .io_out_sum_exp(local_pes_28_21_io_out_sum_exp),
    .io_out_kv(local_pes_28_21_io_out_kv),
    .io_out_stage(local_pes_28_21_io_out_stage)
  );
  PE_1 local_pes_28_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_22_clock),
    .reset(local_pes_28_22_reset),
    .io_in_q(local_pes_28_22_io_in_q),
    .io_in_sum(local_pes_28_22_io_in_sum),
    .io_in_sum_exp(local_pes_28_22_io_in_sum_exp),
    .io_in_kv(local_pes_28_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_22_io_in_inv_sum),
    .io_in_stage(local_pes_28_22_io_in_stage),
    .io_out_q(local_pes_28_22_io_out_q),
    .io_out_sum(local_pes_28_22_io_out_sum),
    .io_out_sum_exp(local_pes_28_22_io_out_sum_exp),
    .io_out_kv(local_pes_28_22_io_out_kv),
    .io_out_stage(local_pes_28_22_io_out_stage)
  );
  PE_1 local_pes_28_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_23_clock),
    .reset(local_pes_28_23_reset),
    .io_in_q(local_pes_28_23_io_in_q),
    .io_in_sum(local_pes_28_23_io_in_sum),
    .io_in_sum_exp(local_pes_28_23_io_in_sum_exp),
    .io_in_kv(local_pes_28_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_23_io_in_inv_sum),
    .io_in_stage(local_pes_28_23_io_in_stage),
    .io_out_q(local_pes_28_23_io_out_q),
    .io_out_sum(local_pes_28_23_io_out_sum),
    .io_out_sum_exp(local_pes_28_23_io_out_sum_exp),
    .io_out_kv(local_pes_28_23_io_out_kv),
    .io_out_stage(local_pes_28_23_io_out_stage)
  );
  PE_1 local_pes_28_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_24_clock),
    .reset(local_pes_28_24_reset),
    .io_in_q(local_pes_28_24_io_in_q),
    .io_in_sum(local_pes_28_24_io_in_sum),
    .io_in_sum_exp(local_pes_28_24_io_in_sum_exp),
    .io_in_kv(local_pes_28_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_24_io_in_inv_sum),
    .io_in_stage(local_pes_28_24_io_in_stage),
    .io_out_q(local_pes_28_24_io_out_q),
    .io_out_sum(local_pes_28_24_io_out_sum),
    .io_out_sum_exp(local_pes_28_24_io_out_sum_exp),
    .io_out_kv(local_pes_28_24_io_out_kv),
    .io_out_stage(local_pes_28_24_io_out_stage)
  );
  PE_1 local_pes_28_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_25_clock),
    .reset(local_pes_28_25_reset),
    .io_in_q(local_pes_28_25_io_in_q),
    .io_in_sum(local_pes_28_25_io_in_sum),
    .io_in_sum_exp(local_pes_28_25_io_in_sum_exp),
    .io_in_kv(local_pes_28_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_25_io_in_inv_sum),
    .io_in_stage(local_pes_28_25_io_in_stage),
    .io_out_q(local_pes_28_25_io_out_q),
    .io_out_sum(local_pes_28_25_io_out_sum),
    .io_out_sum_exp(local_pes_28_25_io_out_sum_exp),
    .io_out_kv(local_pes_28_25_io_out_kv),
    .io_out_stage(local_pes_28_25_io_out_stage)
  );
  PE_1 local_pes_28_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_26_clock),
    .reset(local_pes_28_26_reset),
    .io_in_q(local_pes_28_26_io_in_q),
    .io_in_sum(local_pes_28_26_io_in_sum),
    .io_in_sum_exp(local_pes_28_26_io_in_sum_exp),
    .io_in_kv(local_pes_28_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_26_io_in_inv_sum),
    .io_in_stage(local_pes_28_26_io_in_stage),
    .io_out_q(local_pes_28_26_io_out_q),
    .io_out_sum(local_pes_28_26_io_out_sum),
    .io_out_sum_exp(local_pes_28_26_io_out_sum_exp),
    .io_out_kv(local_pes_28_26_io_out_kv),
    .io_out_stage(local_pes_28_26_io_out_stage)
  );
  PE_1 local_pes_28_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_27_clock),
    .reset(local_pes_28_27_reset),
    .io_in_q(local_pes_28_27_io_in_q),
    .io_in_sum(local_pes_28_27_io_in_sum),
    .io_in_sum_exp(local_pes_28_27_io_in_sum_exp),
    .io_in_kv(local_pes_28_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_27_io_in_inv_sum),
    .io_in_stage(local_pes_28_27_io_in_stage),
    .io_out_q(local_pes_28_27_io_out_q),
    .io_out_sum(local_pes_28_27_io_out_sum),
    .io_out_sum_exp(local_pes_28_27_io_out_sum_exp),
    .io_out_kv(local_pes_28_27_io_out_kv),
    .io_out_stage(local_pes_28_27_io_out_stage)
  );
  PE_1 local_pes_28_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_28_clock),
    .reset(local_pes_28_28_reset),
    .io_in_q(local_pes_28_28_io_in_q),
    .io_in_sum(local_pes_28_28_io_in_sum),
    .io_in_sum_exp(local_pes_28_28_io_in_sum_exp),
    .io_in_kv(local_pes_28_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_28_io_in_inv_sum),
    .io_in_stage(local_pes_28_28_io_in_stage),
    .io_out_q(local_pes_28_28_io_out_q),
    .io_out_sum(local_pes_28_28_io_out_sum),
    .io_out_sum_exp(local_pes_28_28_io_out_sum_exp),
    .io_out_kv(local_pes_28_28_io_out_kv),
    .io_out_stage(local_pes_28_28_io_out_stage)
  );
  PE_1 local_pes_28_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_29_clock),
    .reset(local_pes_28_29_reset),
    .io_in_q(local_pes_28_29_io_in_q),
    .io_in_sum(local_pes_28_29_io_in_sum),
    .io_in_sum_exp(local_pes_28_29_io_in_sum_exp),
    .io_in_kv(local_pes_28_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_29_io_in_inv_sum),
    .io_in_stage(local_pes_28_29_io_in_stage),
    .io_out_q(local_pes_28_29_io_out_q),
    .io_out_sum(local_pes_28_29_io_out_sum),
    .io_out_sum_exp(local_pes_28_29_io_out_sum_exp),
    .io_out_kv(local_pes_28_29_io_out_kv),
    .io_out_stage(local_pes_28_29_io_out_stage)
  );
  PE_1 local_pes_28_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_30_clock),
    .reset(local_pes_28_30_reset),
    .io_in_q(local_pes_28_30_io_in_q),
    .io_in_sum(local_pes_28_30_io_in_sum),
    .io_in_sum_exp(local_pes_28_30_io_in_sum_exp),
    .io_in_kv(local_pes_28_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_30_io_in_inv_sum),
    .io_in_stage(local_pes_28_30_io_in_stage),
    .io_out_q(local_pes_28_30_io_out_q),
    .io_out_sum(local_pes_28_30_io_out_sum),
    .io_out_sum_exp(local_pes_28_30_io_out_sum_exp),
    .io_out_kv(local_pes_28_30_io_out_kv),
    .io_out_stage(local_pes_28_30_io_out_stage)
  );
  PE_1 local_pes_28_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_28_31_clock),
    .reset(local_pes_28_31_reset),
    .io_in_q(local_pes_28_31_io_in_q),
    .io_in_sum(local_pes_28_31_io_in_sum),
    .io_in_sum_exp(local_pes_28_31_io_in_sum_exp),
    .io_in_kv(local_pes_28_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_28_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_28_31_io_in_inv_sum),
    .io_in_stage(local_pes_28_31_io_in_stage),
    .io_out_q(local_pes_28_31_io_out_q),
    .io_out_sum(local_pes_28_31_io_out_sum),
    .io_out_sum_exp(local_pes_28_31_io_out_sum_exp),
    .io_out_kv(local_pes_28_31_io_out_kv),
    .io_out_stage(local_pes_28_31_io_out_stage)
  );
  PE local_pes_29_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_0_clock),
    .reset(local_pes_29_0_reset),
    .io_in_q(local_pes_29_0_io_in_q),
    .io_in_kv(local_pes_29_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_0_io_in_inv_sum),
    .io_in_stage(local_pes_29_0_io_in_stage),
    .io_out_q(local_pes_29_0_io_out_q),
    .io_out_sum(local_pes_29_0_io_out_sum),
    .io_out_kv(local_pes_29_0_io_out_kv),
    .io_out_stage(local_pes_29_0_io_out_stage)
  );
  PE_1 local_pes_29_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_1_clock),
    .reset(local_pes_29_1_reset),
    .io_in_q(local_pes_29_1_io_in_q),
    .io_in_sum(local_pes_29_1_io_in_sum),
    .io_in_sum_exp(local_pes_29_1_io_in_sum_exp),
    .io_in_kv(local_pes_29_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_1_io_in_inv_sum),
    .io_in_stage(local_pes_29_1_io_in_stage),
    .io_out_q(local_pes_29_1_io_out_q),
    .io_out_sum(local_pes_29_1_io_out_sum),
    .io_out_sum_exp(local_pes_29_1_io_out_sum_exp),
    .io_out_kv(local_pes_29_1_io_out_kv),
    .io_out_stage(local_pes_29_1_io_out_stage)
  );
  PE_1 local_pes_29_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_2_clock),
    .reset(local_pes_29_2_reset),
    .io_in_q(local_pes_29_2_io_in_q),
    .io_in_sum(local_pes_29_2_io_in_sum),
    .io_in_sum_exp(local_pes_29_2_io_in_sum_exp),
    .io_in_kv(local_pes_29_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_2_io_in_inv_sum),
    .io_in_stage(local_pes_29_2_io_in_stage),
    .io_out_q(local_pes_29_2_io_out_q),
    .io_out_sum(local_pes_29_2_io_out_sum),
    .io_out_sum_exp(local_pes_29_2_io_out_sum_exp),
    .io_out_kv(local_pes_29_2_io_out_kv),
    .io_out_stage(local_pes_29_2_io_out_stage)
  );
  PE_1 local_pes_29_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_3_clock),
    .reset(local_pes_29_3_reset),
    .io_in_q(local_pes_29_3_io_in_q),
    .io_in_sum(local_pes_29_3_io_in_sum),
    .io_in_sum_exp(local_pes_29_3_io_in_sum_exp),
    .io_in_kv(local_pes_29_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_3_io_in_inv_sum),
    .io_in_stage(local_pes_29_3_io_in_stage),
    .io_out_q(local_pes_29_3_io_out_q),
    .io_out_sum(local_pes_29_3_io_out_sum),
    .io_out_sum_exp(local_pes_29_3_io_out_sum_exp),
    .io_out_kv(local_pes_29_3_io_out_kv),
    .io_out_stage(local_pes_29_3_io_out_stage)
  );
  PE_1 local_pes_29_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_4_clock),
    .reset(local_pes_29_4_reset),
    .io_in_q(local_pes_29_4_io_in_q),
    .io_in_sum(local_pes_29_4_io_in_sum),
    .io_in_sum_exp(local_pes_29_4_io_in_sum_exp),
    .io_in_kv(local_pes_29_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_4_io_in_inv_sum),
    .io_in_stage(local_pes_29_4_io_in_stage),
    .io_out_q(local_pes_29_4_io_out_q),
    .io_out_sum(local_pes_29_4_io_out_sum),
    .io_out_sum_exp(local_pes_29_4_io_out_sum_exp),
    .io_out_kv(local_pes_29_4_io_out_kv),
    .io_out_stage(local_pes_29_4_io_out_stage)
  );
  PE_1 local_pes_29_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_5_clock),
    .reset(local_pes_29_5_reset),
    .io_in_q(local_pes_29_5_io_in_q),
    .io_in_sum(local_pes_29_5_io_in_sum),
    .io_in_sum_exp(local_pes_29_5_io_in_sum_exp),
    .io_in_kv(local_pes_29_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_5_io_in_inv_sum),
    .io_in_stage(local_pes_29_5_io_in_stage),
    .io_out_q(local_pes_29_5_io_out_q),
    .io_out_sum(local_pes_29_5_io_out_sum),
    .io_out_sum_exp(local_pes_29_5_io_out_sum_exp),
    .io_out_kv(local_pes_29_5_io_out_kv),
    .io_out_stage(local_pes_29_5_io_out_stage)
  );
  PE_1 local_pes_29_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_6_clock),
    .reset(local_pes_29_6_reset),
    .io_in_q(local_pes_29_6_io_in_q),
    .io_in_sum(local_pes_29_6_io_in_sum),
    .io_in_sum_exp(local_pes_29_6_io_in_sum_exp),
    .io_in_kv(local_pes_29_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_6_io_in_inv_sum),
    .io_in_stage(local_pes_29_6_io_in_stage),
    .io_out_q(local_pes_29_6_io_out_q),
    .io_out_sum(local_pes_29_6_io_out_sum),
    .io_out_sum_exp(local_pes_29_6_io_out_sum_exp),
    .io_out_kv(local_pes_29_6_io_out_kv),
    .io_out_stage(local_pes_29_6_io_out_stage)
  );
  PE_1 local_pes_29_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_7_clock),
    .reset(local_pes_29_7_reset),
    .io_in_q(local_pes_29_7_io_in_q),
    .io_in_sum(local_pes_29_7_io_in_sum),
    .io_in_sum_exp(local_pes_29_7_io_in_sum_exp),
    .io_in_kv(local_pes_29_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_7_io_in_inv_sum),
    .io_in_stage(local_pes_29_7_io_in_stage),
    .io_out_q(local_pes_29_7_io_out_q),
    .io_out_sum(local_pes_29_7_io_out_sum),
    .io_out_sum_exp(local_pes_29_7_io_out_sum_exp),
    .io_out_kv(local_pes_29_7_io_out_kv),
    .io_out_stage(local_pes_29_7_io_out_stage)
  );
  PE_1 local_pes_29_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_8_clock),
    .reset(local_pes_29_8_reset),
    .io_in_q(local_pes_29_8_io_in_q),
    .io_in_sum(local_pes_29_8_io_in_sum),
    .io_in_sum_exp(local_pes_29_8_io_in_sum_exp),
    .io_in_kv(local_pes_29_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_8_io_in_inv_sum),
    .io_in_stage(local_pes_29_8_io_in_stage),
    .io_out_q(local_pes_29_8_io_out_q),
    .io_out_sum(local_pes_29_8_io_out_sum),
    .io_out_sum_exp(local_pes_29_8_io_out_sum_exp),
    .io_out_kv(local_pes_29_8_io_out_kv),
    .io_out_stage(local_pes_29_8_io_out_stage)
  );
  PE_1 local_pes_29_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_9_clock),
    .reset(local_pes_29_9_reset),
    .io_in_q(local_pes_29_9_io_in_q),
    .io_in_sum(local_pes_29_9_io_in_sum),
    .io_in_sum_exp(local_pes_29_9_io_in_sum_exp),
    .io_in_kv(local_pes_29_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_9_io_in_inv_sum),
    .io_in_stage(local_pes_29_9_io_in_stage),
    .io_out_q(local_pes_29_9_io_out_q),
    .io_out_sum(local_pes_29_9_io_out_sum),
    .io_out_sum_exp(local_pes_29_9_io_out_sum_exp),
    .io_out_kv(local_pes_29_9_io_out_kv),
    .io_out_stage(local_pes_29_9_io_out_stage)
  );
  PE_1 local_pes_29_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_10_clock),
    .reset(local_pes_29_10_reset),
    .io_in_q(local_pes_29_10_io_in_q),
    .io_in_sum(local_pes_29_10_io_in_sum),
    .io_in_sum_exp(local_pes_29_10_io_in_sum_exp),
    .io_in_kv(local_pes_29_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_10_io_in_inv_sum),
    .io_in_stage(local_pes_29_10_io_in_stage),
    .io_out_q(local_pes_29_10_io_out_q),
    .io_out_sum(local_pes_29_10_io_out_sum),
    .io_out_sum_exp(local_pes_29_10_io_out_sum_exp),
    .io_out_kv(local_pes_29_10_io_out_kv),
    .io_out_stage(local_pes_29_10_io_out_stage)
  );
  PE_1 local_pes_29_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_11_clock),
    .reset(local_pes_29_11_reset),
    .io_in_q(local_pes_29_11_io_in_q),
    .io_in_sum(local_pes_29_11_io_in_sum),
    .io_in_sum_exp(local_pes_29_11_io_in_sum_exp),
    .io_in_kv(local_pes_29_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_11_io_in_inv_sum),
    .io_in_stage(local_pes_29_11_io_in_stage),
    .io_out_q(local_pes_29_11_io_out_q),
    .io_out_sum(local_pes_29_11_io_out_sum),
    .io_out_sum_exp(local_pes_29_11_io_out_sum_exp),
    .io_out_kv(local_pes_29_11_io_out_kv),
    .io_out_stage(local_pes_29_11_io_out_stage)
  );
  PE_1 local_pes_29_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_12_clock),
    .reset(local_pes_29_12_reset),
    .io_in_q(local_pes_29_12_io_in_q),
    .io_in_sum(local_pes_29_12_io_in_sum),
    .io_in_sum_exp(local_pes_29_12_io_in_sum_exp),
    .io_in_kv(local_pes_29_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_12_io_in_inv_sum),
    .io_in_stage(local_pes_29_12_io_in_stage),
    .io_out_q(local_pes_29_12_io_out_q),
    .io_out_sum(local_pes_29_12_io_out_sum),
    .io_out_sum_exp(local_pes_29_12_io_out_sum_exp),
    .io_out_kv(local_pes_29_12_io_out_kv),
    .io_out_stage(local_pes_29_12_io_out_stage)
  );
  PE_1 local_pes_29_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_13_clock),
    .reset(local_pes_29_13_reset),
    .io_in_q(local_pes_29_13_io_in_q),
    .io_in_sum(local_pes_29_13_io_in_sum),
    .io_in_sum_exp(local_pes_29_13_io_in_sum_exp),
    .io_in_kv(local_pes_29_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_13_io_in_inv_sum),
    .io_in_stage(local_pes_29_13_io_in_stage),
    .io_out_q(local_pes_29_13_io_out_q),
    .io_out_sum(local_pes_29_13_io_out_sum),
    .io_out_sum_exp(local_pes_29_13_io_out_sum_exp),
    .io_out_kv(local_pes_29_13_io_out_kv),
    .io_out_stage(local_pes_29_13_io_out_stage)
  );
  PE_1 local_pes_29_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_14_clock),
    .reset(local_pes_29_14_reset),
    .io_in_q(local_pes_29_14_io_in_q),
    .io_in_sum(local_pes_29_14_io_in_sum),
    .io_in_sum_exp(local_pes_29_14_io_in_sum_exp),
    .io_in_kv(local_pes_29_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_14_io_in_inv_sum),
    .io_in_stage(local_pes_29_14_io_in_stage),
    .io_out_q(local_pes_29_14_io_out_q),
    .io_out_sum(local_pes_29_14_io_out_sum),
    .io_out_sum_exp(local_pes_29_14_io_out_sum_exp),
    .io_out_kv(local_pes_29_14_io_out_kv),
    .io_out_stage(local_pes_29_14_io_out_stage)
  );
  PE_1 local_pes_29_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_15_clock),
    .reset(local_pes_29_15_reset),
    .io_in_q(local_pes_29_15_io_in_q),
    .io_in_sum(local_pes_29_15_io_in_sum),
    .io_in_sum_exp(local_pes_29_15_io_in_sum_exp),
    .io_in_kv(local_pes_29_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_15_io_in_inv_sum),
    .io_in_stage(local_pes_29_15_io_in_stage),
    .io_out_q(local_pes_29_15_io_out_q),
    .io_out_sum(local_pes_29_15_io_out_sum),
    .io_out_sum_exp(local_pes_29_15_io_out_sum_exp),
    .io_out_kv(local_pes_29_15_io_out_kv),
    .io_out_stage(local_pes_29_15_io_out_stage)
  );
  PE_1 local_pes_29_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_16_clock),
    .reset(local_pes_29_16_reset),
    .io_in_q(local_pes_29_16_io_in_q),
    .io_in_sum(local_pes_29_16_io_in_sum),
    .io_in_sum_exp(local_pes_29_16_io_in_sum_exp),
    .io_in_kv(local_pes_29_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_16_io_in_inv_sum),
    .io_in_stage(local_pes_29_16_io_in_stage),
    .io_out_q(local_pes_29_16_io_out_q),
    .io_out_sum(local_pes_29_16_io_out_sum),
    .io_out_sum_exp(local_pes_29_16_io_out_sum_exp),
    .io_out_kv(local_pes_29_16_io_out_kv),
    .io_out_stage(local_pes_29_16_io_out_stage)
  );
  PE_1 local_pes_29_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_17_clock),
    .reset(local_pes_29_17_reset),
    .io_in_q(local_pes_29_17_io_in_q),
    .io_in_sum(local_pes_29_17_io_in_sum),
    .io_in_sum_exp(local_pes_29_17_io_in_sum_exp),
    .io_in_kv(local_pes_29_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_17_io_in_inv_sum),
    .io_in_stage(local_pes_29_17_io_in_stage),
    .io_out_q(local_pes_29_17_io_out_q),
    .io_out_sum(local_pes_29_17_io_out_sum),
    .io_out_sum_exp(local_pes_29_17_io_out_sum_exp),
    .io_out_kv(local_pes_29_17_io_out_kv),
    .io_out_stage(local_pes_29_17_io_out_stage)
  );
  PE_1 local_pes_29_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_18_clock),
    .reset(local_pes_29_18_reset),
    .io_in_q(local_pes_29_18_io_in_q),
    .io_in_sum(local_pes_29_18_io_in_sum),
    .io_in_sum_exp(local_pes_29_18_io_in_sum_exp),
    .io_in_kv(local_pes_29_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_18_io_in_inv_sum),
    .io_in_stage(local_pes_29_18_io_in_stage),
    .io_out_q(local_pes_29_18_io_out_q),
    .io_out_sum(local_pes_29_18_io_out_sum),
    .io_out_sum_exp(local_pes_29_18_io_out_sum_exp),
    .io_out_kv(local_pes_29_18_io_out_kv),
    .io_out_stage(local_pes_29_18_io_out_stage)
  );
  PE_1 local_pes_29_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_19_clock),
    .reset(local_pes_29_19_reset),
    .io_in_q(local_pes_29_19_io_in_q),
    .io_in_sum(local_pes_29_19_io_in_sum),
    .io_in_sum_exp(local_pes_29_19_io_in_sum_exp),
    .io_in_kv(local_pes_29_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_19_io_in_inv_sum),
    .io_in_stage(local_pes_29_19_io_in_stage),
    .io_out_q(local_pes_29_19_io_out_q),
    .io_out_sum(local_pes_29_19_io_out_sum),
    .io_out_sum_exp(local_pes_29_19_io_out_sum_exp),
    .io_out_kv(local_pes_29_19_io_out_kv),
    .io_out_stage(local_pes_29_19_io_out_stage)
  );
  PE_1 local_pes_29_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_20_clock),
    .reset(local_pes_29_20_reset),
    .io_in_q(local_pes_29_20_io_in_q),
    .io_in_sum(local_pes_29_20_io_in_sum),
    .io_in_sum_exp(local_pes_29_20_io_in_sum_exp),
    .io_in_kv(local_pes_29_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_20_io_in_inv_sum),
    .io_in_stage(local_pes_29_20_io_in_stage),
    .io_out_q(local_pes_29_20_io_out_q),
    .io_out_sum(local_pes_29_20_io_out_sum),
    .io_out_sum_exp(local_pes_29_20_io_out_sum_exp),
    .io_out_kv(local_pes_29_20_io_out_kv),
    .io_out_stage(local_pes_29_20_io_out_stage)
  );
  PE_1 local_pes_29_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_21_clock),
    .reset(local_pes_29_21_reset),
    .io_in_q(local_pes_29_21_io_in_q),
    .io_in_sum(local_pes_29_21_io_in_sum),
    .io_in_sum_exp(local_pes_29_21_io_in_sum_exp),
    .io_in_kv(local_pes_29_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_21_io_in_inv_sum),
    .io_in_stage(local_pes_29_21_io_in_stage),
    .io_out_q(local_pes_29_21_io_out_q),
    .io_out_sum(local_pes_29_21_io_out_sum),
    .io_out_sum_exp(local_pes_29_21_io_out_sum_exp),
    .io_out_kv(local_pes_29_21_io_out_kv),
    .io_out_stage(local_pes_29_21_io_out_stage)
  );
  PE_1 local_pes_29_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_22_clock),
    .reset(local_pes_29_22_reset),
    .io_in_q(local_pes_29_22_io_in_q),
    .io_in_sum(local_pes_29_22_io_in_sum),
    .io_in_sum_exp(local_pes_29_22_io_in_sum_exp),
    .io_in_kv(local_pes_29_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_22_io_in_inv_sum),
    .io_in_stage(local_pes_29_22_io_in_stage),
    .io_out_q(local_pes_29_22_io_out_q),
    .io_out_sum(local_pes_29_22_io_out_sum),
    .io_out_sum_exp(local_pes_29_22_io_out_sum_exp),
    .io_out_kv(local_pes_29_22_io_out_kv),
    .io_out_stage(local_pes_29_22_io_out_stage)
  );
  PE_1 local_pes_29_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_23_clock),
    .reset(local_pes_29_23_reset),
    .io_in_q(local_pes_29_23_io_in_q),
    .io_in_sum(local_pes_29_23_io_in_sum),
    .io_in_sum_exp(local_pes_29_23_io_in_sum_exp),
    .io_in_kv(local_pes_29_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_23_io_in_inv_sum),
    .io_in_stage(local_pes_29_23_io_in_stage),
    .io_out_q(local_pes_29_23_io_out_q),
    .io_out_sum(local_pes_29_23_io_out_sum),
    .io_out_sum_exp(local_pes_29_23_io_out_sum_exp),
    .io_out_kv(local_pes_29_23_io_out_kv),
    .io_out_stage(local_pes_29_23_io_out_stage)
  );
  PE_1 local_pes_29_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_24_clock),
    .reset(local_pes_29_24_reset),
    .io_in_q(local_pes_29_24_io_in_q),
    .io_in_sum(local_pes_29_24_io_in_sum),
    .io_in_sum_exp(local_pes_29_24_io_in_sum_exp),
    .io_in_kv(local_pes_29_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_24_io_in_inv_sum),
    .io_in_stage(local_pes_29_24_io_in_stage),
    .io_out_q(local_pes_29_24_io_out_q),
    .io_out_sum(local_pes_29_24_io_out_sum),
    .io_out_sum_exp(local_pes_29_24_io_out_sum_exp),
    .io_out_kv(local_pes_29_24_io_out_kv),
    .io_out_stage(local_pes_29_24_io_out_stage)
  );
  PE_1 local_pes_29_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_25_clock),
    .reset(local_pes_29_25_reset),
    .io_in_q(local_pes_29_25_io_in_q),
    .io_in_sum(local_pes_29_25_io_in_sum),
    .io_in_sum_exp(local_pes_29_25_io_in_sum_exp),
    .io_in_kv(local_pes_29_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_25_io_in_inv_sum),
    .io_in_stage(local_pes_29_25_io_in_stage),
    .io_out_q(local_pes_29_25_io_out_q),
    .io_out_sum(local_pes_29_25_io_out_sum),
    .io_out_sum_exp(local_pes_29_25_io_out_sum_exp),
    .io_out_kv(local_pes_29_25_io_out_kv),
    .io_out_stage(local_pes_29_25_io_out_stage)
  );
  PE_1 local_pes_29_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_26_clock),
    .reset(local_pes_29_26_reset),
    .io_in_q(local_pes_29_26_io_in_q),
    .io_in_sum(local_pes_29_26_io_in_sum),
    .io_in_sum_exp(local_pes_29_26_io_in_sum_exp),
    .io_in_kv(local_pes_29_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_26_io_in_inv_sum),
    .io_in_stage(local_pes_29_26_io_in_stage),
    .io_out_q(local_pes_29_26_io_out_q),
    .io_out_sum(local_pes_29_26_io_out_sum),
    .io_out_sum_exp(local_pes_29_26_io_out_sum_exp),
    .io_out_kv(local_pes_29_26_io_out_kv),
    .io_out_stage(local_pes_29_26_io_out_stage)
  );
  PE_1 local_pes_29_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_27_clock),
    .reset(local_pes_29_27_reset),
    .io_in_q(local_pes_29_27_io_in_q),
    .io_in_sum(local_pes_29_27_io_in_sum),
    .io_in_sum_exp(local_pes_29_27_io_in_sum_exp),
    .io_in_kv(local_pes_29_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_27_io_in_inv_sum),
    .io_in_stage(local_pes_29_27_io_in_stage),
    .io_out_q(local_pes_29_27_io_out_q),
    .io_out_sum(local_pes_29_27_io_out_sum),
    .io_out_sum_exp(local_pes_29_27_io_out_sum_exp),
    .io_out_kv(local_pes_29_27_io_out_kv),
    .io_out_stage(local_pes_29_27_io_out_stage)
  );
  PE_1 local_pes_29_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_28_clock),
    .reset(local_pes_29_28_reset),
    .io_in_q(local_pes_29_28_io_in_q),
    .io_in_sum(local_pes_29_28_io_in_sum),
    .io_in_sum_exp(local_pes_29_28_io_in_sum_exp),
    .io_in_kv(local_pes_29_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_28_io_in_inv_sum),
    .io_in_stage(local_pes_29_28_io_in_stage),
    .io_out_q(local_pes_29_28_io_out_q),
    .io_out_sum(local_pes_29_28_io_out_sum),
    .io_out_sum_exp(local_pes_29_28_io_out_sum_exp),
    .io_out_kv(local_pes_29_28_io_out_kv),
    .io_out_stage(local_pes_29_28_io_out_stage)
  );
  PE_1 local_pes_29_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_29_clock),
    .reset(local_pes_29_29_reset),
    .io_in_q(local_pes_29_29_io_in_q),
    .io_in_sum(local_pes_29_29_io_in_sum),
    .io_in_sum_exp(local_pes_29_29_io_in_sum_exp),
    .io_in_kv(local_pes_29_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_29_io_in_inv_sum),
    .io_in_stage(local_pes_29_29_io_in_stage),
    .io_out_q(local_pes_29_29_io_out_q),
    .io_out_sum(local_pes_29_29_io_out_sum),
    .io_out_sum_exp(local_pes_29_29_io_out_sum_exp),
    .io_out_kv(local_pes_29_29_io_out_kv),
    .io_out_stage(local_pes_29_29_io_out_stage)
  );
  PE_1 local_pes_29_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_30_clock),
    .reset(local_pes_29_30_reset),
    .io_in_q(local_pes_29_30_io_in_q),
    .io_in_sum(local_pes_29_30_io_in_sum),
    .io_in_sum_exp(local_pes_29_30_io_in_sum_exp),
    .io_in_kv(local_pes_29_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_30_io_in_inv_sum),
    .io_in_stage(local_pes_29_30_io_in_stage),
    .io_out_q(local_pes_29_30_io_out_q),
    .io_out_sum(local_pes_29_30_io_out_sum),
    .io_out_sum_exp(local_pes_29_30_io_out_sum_exp),
    .io_out_kv(local_pes_29_30_io_out_kv),
    .io_out_stage(local_pes_29_30_io_out_stage)
  );
  PE_1 local_pes_29_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_29_31_clock),
    .reset(local_pes_29_31_reset),
    .io_in_q(local_pes_29_31_io_in_q),
    .io_in_sum(local_pes_29_31_io_in_sum),
    .io_in_sum_exp(local_pes_29_31_io_in_sum_exp),
    .io_in_kv(local_pes_29_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_29_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_29_31_io_in_inv_sum),
    .io_in_stage(local_pes_29_31_io_in_stage),
    .io_out_q(local_pes_29_31_io_out_q),
    .io_out_sum(local_pes_29_31_io_out_sum),
    .io_out_sum_exp(local_pes_29_31_io_out_sum_exp),
    .io_out_kv(local_pes_29_31_io_out_kv),
    .io_out_stage(local_pes_29_31_io_out_stage)
  );
  PE local_pes_30_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_0_clock),
    .reset(local_pes_30_0_reset),
    .io_in_q(local_pes_30_0_io_in_q),
    .io_in_kv(local_pes_30_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_0_io_in_inv_sum),
    .io_in_stage(local_pes_30_0_io_in_stage),
    .io_out_q(local_pes_30_0_io_out_q),
    .io_out_sum(local_pes_30_0_io_out_sum),
    .io_out_kv(local_pes_30_0_io_out_kv),
    .io_out_stage(local_pes_30_0_io_out_stage)
  );
  PE_1 local_pes_30_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_1_clock),
    .reset(local_pes_30_1_reset),
    .io_in_q(local_pes_30_1_io_in_q),
    .io_in_sum(local_pes_30_1_io_in_sum),
    .io_in_sum_exp(local_pes_30_1_io_in_sum_exp),
    .io_in_kv(local_pes_30_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_1_io_in_inv_sum),
    .io_in_stage(local_pes_30_1_io_in_stage),
    .io_out_q(local_pes_30_1_io_out_q),
    .io_out_sum(local_pes_30_1_io_out_sum),
    .io_out_sum_exp(local_pes_30_1_io_out_sum_exp),
    .io_out_kv(local_pes_30_1_io_out_kv),
    .io_out_stage(local_pes_30_1_io_out_stage)
  );
  PE_1 local_pes_30_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_2_clock),
    .reset(local_pes_30_2_reset),
    .io_in_q(local_pes_30_2_io_in_q),
    .io_in_sum(local_pes_30_2_io_in_sum),
    .io_in_sum_exp(local_pes_30_2_io_in_sum_exp),
    .io_in_kv(local_pes_30_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_2_io_in_inv_sum),
    .io_in_stage(local_pes_30_2_io_in_stage),
    .io_out_q(local_pes_30_2_io_out_q),
    .io_out_sum(local_pes_30_2_io_out_sum),
    .io_out_sum_exp(local_pes_30_2_io_out_sum_exp),
    .io_out_kv(local_pes_30_2_io_out_kv),
    .io_out_stage(local_pes_30_2_io_out_stage)
  );
  PE_1 local_pes_30_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_3_clock),
    .reset(local_pes_30_3_reset),
    .io_in_q(local_pes_30_3_io_in_q),
    .io_in_sum(local_pes_30_3_io_in_sum),
    .io_in_sum_exp(local_pes_30_3_io_in_sum_exp),
    .io_in_kv(local_pes_30_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_3_io_in_inv_sum),
    .io_in_stage(local_pes_30_3_io_in_stage),
    .io_out_q(local_pes_30_3_io_out_q),
    .io_out_sum(local_pes_30_3_io_out_sum),
    .io_out_sum_exp(local_pes_30_3_io_out_sum_exp),
    .io_out_kv(local_pes_30_3_io_out_kv),
    .io_out_stage(local_pes_30_3_io_out_stage)
  );
  PE_1 local_pes_30_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_4_clock),
    .reset(local_pes_30_4_reset),
    .io_in_q(local_pes_30_4_io_in_q),
    .io_in_sum(local_pes_30_4_io_in_sum),
    .io_in_sum_exp(local_pes_30_4_io_in_sum_exp),
    .io_in_kv(local_pes_30_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_4_io_in_inv_sum),
    .io_in_stage(local_pes_30_4_io_in_stage),
    .io_out_q(local_pes_30_4_io_out_q),
    .io_out_sum(local_pes_30_4_io_out_sum),
    .io_out_sum_exp(local_pes_30_4_io_out_sum_exp),
    .io_out_kv(local_pes_30_4_io_out_kv),
    .io_out_stage(local_pes_30_4_io_out_stage)
  );
  PE_1 local_pes_30_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_5_clock),
    .reset(local_pes_30_5_reset),
    .io_in_q(local_pes_30_5_io_in_q),
    .io_in_sum(local_pes_30_5_io_in_sum),
    .io_in_sum_exp(local_pes_30_5_io_in_sum_exp),
    .io_in_kv(local_pes_30_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_5_io_in_inv_sum),
    .io_in_stage(local_pes_30_5_io_in_stage),
    .io_out_q(local_pes_30_5_io_out_q),
    .io_out_sum(local_pes_30_5_io_out_sum),
    .io_out_sum_exp(local_pes_30_5_io_out_sum_exp),
    .io_out_kv(local_pes_30_5_io_out_kv),
    .io_out_stage(local_pes_30_5_io_out_stage)
  );
  PE_1 local_pes_30_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_6_clock),
    .reset(local_pes_30_6_reset),
    .io_in_q(local_pes_30_6_io_in_q),
    .io_in_sum(local_pes_30_6_io_in_sum),
    .io_in_sum_exp(local_pes_30_6_io_in_sum_exp),
    .io_in_kv(local_pes_30_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_6_io_in_inv_sum),
    .io_in_stage(local_pes_30_6_io_in_stage),
    .io_out_q(local_pes_30_6_io_out_q),
    .io_out_sum(local_pes_30_6_io_out_sum),
    .io_out_sum_exp(local_pes_30_6_io_out_sum_exp),
    .io_out_kv(local_pes_30_6_io_out_kv),
    .io_out_stage(local_pes_30_6_io_out_stage)
  );
  PE_1 local_pes_30_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_7_clock),
    .reset(local_pes_30_7_reset),
    .io_in_q(local_pes_30_7_io_in_q),
    .io_in_sum(local_pes_30_7_io_in_sum),
    .io_in_sum_exp(local_pes_30_7_io_in_sum_exp),
    .io_in_kv(local_pes_30_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_7_io_in_inv_sum),
    .io_in_stage(local_pes_30_7_io_in_stage),
    .io_out_q(local_pes_30_7_io_out_q),
    .io_out_sum(local_pes_30_7_io_out_sum),
    .io_out_sum_exp(local_pes_30_7_io_out_sum_exp),
    .io_out_kv(local_pes_30_7_io_out_kv),
    .io_out_stage(local_pes_30_7_io_out_stage)
  );
  PE_1 local_pes_30_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_8_clock),
    .reset(local_pes_30_8_reset),
    .io_in_q(local_pes_30_8_io_in_q),
    .io_in_sum(local_pes_30_8_io_in_sum),
    .io_in_sum_exp(local_pes_30_8_io_in_sum_exp),
    .io_in_kv(local_pes_30_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_8_io_in_inv_sum),
    .io_in_stage(local_pes_30_8_io_in_stage),
    .io_out_q(local_pes_30_8_io_out_q),
    .io_out_sum(local_pes_30_8_io_out_sum),
    .io_out_sum_exp(local_pes_30_8_io_out_sum_exp),
    .io_out_kv(local_pes_30_8_io_out_kv),
    .io_out_stage(local_pes_30_8_io_out_stage)
  );
  PE_1 local_pes_30_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_9_clock),
    .reset(local_pes_30_9_reset),
    .io_in_q(local_pes_30_9_io_in_q),
    .io_in_sum(local_pes_30_9_io_in_sum),
    .io_in_sum_exp(local_pes_30_9_io_in_sum_exp),
    .io_in_kv(local_pes_30_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_9_io_in_inv_sum),
    .io_in_stage(local_pes_30_9_io_in_stage),
    .io_out_q(local_pes_30_9_io_out_q),
    .io_out_sum(local_pes_30_9_io_out_sum),
    .io_out_sum_exp(local_pes_30_9_io_out_sum_exp),
    .io_out_kv(local_pes_30_9_io_out_kv),
    .io_out_stage(local_pes_30_9_io_out_stage)
  );
  PE_1 local_pes_30_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_10_clock),
    .reset(local_pes_30_10_reset),
    .io_in_q(local_pes_30_10_io_in_q),
    .io_in_sum(local_pes_30_10_io_in_sum),
    .io_in_sum_exp(local_pes_30_10_io_in_sum_exp),
    .io_in_kv(local_pes_30_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_10_io_in_inv_sum),
    .io_in_stage(local_pes_30_10_io_in_stage),
    .io_out_q(local_pes_30_10_io_out_q),
    .io_out_sum(local_pes_30_10_io_out_sum),
    .io_out_sum_exp(local_pes_30_10_io_out_sum_exp),
    .io_out_kv(local_pes_30_10_io_out_kv),
    .io_out_stage(local_pes_30_10_io_out_stage)
  );
  PE_1 local_pes_30_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_11_clock),
    .reset(local_pes_30_11_reset),
    .io_in_q(local_pes_30_11_io_in_q),
    .io_in_sum(local_pes_30_11_io_in_sum),
    .io_in_sum_exp(local_pes_30_11_io_in_sum_exp),
    .io_in_kv(local_pes_30_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_11_io_in_inv_sum),
    .io_in_stage(local_pes_30_11_io_in_stage),
    .io_out_q(local_pes_30_11_io_out_q),
    .io_out_sum(local_pes_30_11_io_out_sum),
    .io_out_sum_exp(local_pes_30_11_io_out_sum_exp),
    .io_out_kv(local_pes_30_11_io_out_kv),
    .io_out_stage(local_pes_30_11_io_out_stage)
  );
  PE_1 local_pes_30_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_12_clock),
    .reset(local_pes_30_12_reset),
    .io_in_q(local_pes_30_12_io_in_q),
    .io_in_sum(local_pes_30_12_io_in_sum),
    .io_in_sum_exp(local_pes_30_12_io_in_sum_exp),
    .io_in_kv(local_pes_30_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_12_io_in_inv_sum),
    .io_in_stage(local_pes_30_12_io_in_stage),
    .io_out_q(local_pes_30_12_io_out_q),
    .io_out_sum(local_pes_30_12_io_out_sum),
    .io_out_sum_exp(local_pes_30_12_io_out_sum_exp),
    .io_out_kv(local_pes_30_12_io_out_kv),
    .io_out_stage(local_pes_30_12_io_out_stage)
  );
  PE_1 local_pes_30_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_13_clock),
    .reset(local_pes_30_13_reset),
    .io_in_q(local_pes_30_13_io_in_q),
    .io_in_sum(local_pes_30_13_io_in_sum),
    .io_in_sum_exp(local_pes_30_13_io_in_sum_exp),
    .io_in_kv(local_pes_30_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_13_io_in_inv_sum),
    .io_in_stage(local_pes_30_13_io_in_stage),
    .io_out_q(local_pes_30_13_io_out_q),
    .io_out_sum(local_pes_30_13_io_out_sum),
    .io_out_sum_exp(local_pes_30_13_io_out_sum_exp),
    .io_out_kv(local_pes_30_13_io_out_kv),
    .io_out_stage(local_pes_30_13_io_out_stage)
  );
  PE_1 local_pes_30_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_14_clock),
    .reset(local_pes_30_14_reset),
    .io_in_q(local_pes_30_14_io_in_q),
    .io_in_sum(local_pes_30_14_io_in_sum),
    .io_in_sum_exp(local_pes_30_14_io_in_sum_exp),
    .io_in_kv(local_pes_30_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_14_io_in_inv_sum),
    .io_in_stage(local_pes_30_14_io_in_stage),
    .io_out_q(local_pes_30_14_io_out_q),
    .io_out_sum(local_pes_30_14_io_out_sum),
    .io_out_sum_exp(local_pes_30_14_io_out_sum_exp),
    .io_out_kv(local_pes_30_14_io_out_kv),
    .io_out_stage(local_pes_30_14_io_out_stage)
  );
  PE_1 local_pes_30_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_15_clock),
    .reset(local_pes_30_15_reset),
    .io_in_q(local_pes_30_15_io_in_q),
    .io_in_sum(local_pes_30_15_io_in_sum),
    .io_in_sum_exp(local_pes_30_15_io_in_sum_exp),
    .io_in_kv(local_pes_30_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_15_io_in_inv_sum),
    .io_in_stage(local_pes_30_15_io_in_stage),
    .io_out_q(local_pes_30_15_io_out_q),
    .io_out_sum(local_pes_30_15_io_out_sum),
    .io_out_sum_exp(local_pes_30_15_io_out_sum_exp),
    .io_out_kv(local_pes_30_15_io_out_kv),
    .io_out_stage(local_pes_30_15_io_out_stage)
  );
  PE_1 local_pes_30_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_16_clock),
    .reset(local_pes_30_16_reset),
    .io_in_q(local_pes_30_16_io_in_q),
    .io_in_sum(local_pes_30_16_io_in_sum),
    .io_in_sum_exp(local_pes_30_16_io_in_sum_exp),
    .io_in_kv(local_pes_30_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_16_io_in_inv_sum),
    .io_in_stage(local_pes_30_16_io_in_stage),
    .io_out_q(local_pes_30_16_io_out_q),
    .io_out_sum(local_pes_30_16_io_out_sum),
    .io_out_sum_exp(local_pes_30_16_io_out_sum_exp),
    .io_out_kv(local_pes_30_16_io_out_kv),
    .io_out_stage(local_pes_30_16_io_out_stage)
  );
  PE_1 local_pes_30_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_17_clock),
    .reset(local_pes_30_17_reset),
    .io_in_q(local_pes_30_17_io_in_q),
    .io_in_sum(local_pes_30_17_io_in_sum),
    .io_in_sum_exp(local_pes_30_17_io_in_sum_exp),
    .io_in_kv(local_pes_30_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_17_io_in_inv_sum),
    .io_in_stage(local_pes_30_17_io_in_stage),
    .io_out_q(local_pes_30_17_io_out_q),
    .io_out_sum(local_pes_30_17_io_out_sum),
    .io_out_sum_exp(local_pes_30_17_io_out_sum_exp),
    .io_out_kv(local_pes_30_17_io_out_kv),
    .io_out_stage(local_pes_30_17_io_out_stage)
  );
  PE_1 local_pes_30_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_18_clock),
    .reset(local_pes_30_18_reset),
    .io_in_q(local_pes_30_18_io_in_q),
    .io_in_sum(local_pes_30_18_io_in_sum),
    .io_in_sum_exp(local_pes_30_18_io_in_sum_exp),
    .io_in_kv(local_pes_30_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_18_io_in_inv_sum),
    .io_in_stage(local_pes_30_18_io_in_stage),
    .io_out_q(local_pes_30_18_io_out_q),
    .io_out_sum(local_pes_30_18_io_out_sum),
    .io_out_sum_exp(local_pes_30_18_io_out_sum_exp),
    .io_out_kv(local_pes_30_18_io_out_kv),
    .io_out_stage(local_pes_30_18_io_out_stage)
  );
  PE_1 local_pes_30_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_19_clock),
    .reset(local_pes_30_19_reset),
    .io_in_q(local_pes_30_19_io_in_q),
    .io_in_sum(local_pes_30_19_io_in_sum),
    .io_in_sum_exp(local_pes_30_19_io_in_sum_exp),
    .io_in_kv(local_pes_30_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_19_io_in_inv_sum),
    .io_in_stage(local_pes_30_19_io_in_stage),
    .io_out_q(local_pes_30_19_io_out_q),
    .io_out_sum(local_pes_30_19_io_out_sum),
    .io_out_sum_exp(local_pes_30_19_io_out_sum_exp),
    .io_out_kv(local_pes_30_19_io_out_kv),
    .io_out_stage(local_pes_30_19_io_out_stage)
  );
  PE_1 local_pes_30_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_20_clock),
    .reset(local_pes_30_20_reset),
    .io_in_q(local_pes_30_20_io_in_q),
    .io_in_sum(local_pes_30_20_io_in_sum),
    .io_in_sum_exp(local_pes_30_20_io_in_sum_exp),
    .io_in_kv(local_pes_30_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_20_io_in_inv_sum),
    .io_in_stage(local_pes_30_20_io_in_stage),
    .io_out_q(local_pes_30_20_io_out_q),
    .io_out_sum(local_pes_30_20_io_out_sum),
    .io_out_sum_exp(local_pes_30_20_io_out_sum_exp),
    .io_out_kv(local_pes_30_20_io_out_kv),
    .io_out_stage(local_pes_30_20_io_out_stage)
  );
  PE_1 local_pes_30_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_21_clock),
    .reset(local_pes_30_21_reset),
    .io_in_q(local_pes_30_21_io_in_q),
    .io_in_sum(local_pes_30_21_io_in_sum),
    .io_in_sum_exp(local_pes_30_21_io_in_sum_exp),
    .io_in_kv(local_pes_30_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_21_io_in_inv_sum),
    .io_in_stage(local_pes_30_21_io_in_stage),
    .io_out_q(local_pes_30_21_io_out_q),
    .io_out_sum(local_pes_30_21_io_out_sum),
    .io_out_sum_exp(local_pes_30_21_io_out_sum_exp),
    .io_out_kv(local_pes_30_21_io_out_kv),
    .io_out_stage(local_pes_30_21_io_out_stage)
  );
  PE_1 local_pes_30_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_22_clock),
    .reset(local_pes_30_22_reset),
    .io_in_q(local_pes_30_22_io_in_q),
    .io_in_sum(local_pes_30_22_io_in_sum),
    .io_in_sum_exp(local_pes_30_22_io_in_sum_exp),
    .io_in_kv(local_pes_30_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_22_io_in_inv_sum),
    .io_in_stage(local_pes_30_22_io_in_stage),
    .io_out_q(local_pes_30_22_io_out_q),
    .io_out_sum(local_pes_30_22_io_out_sum),
    .io_out_sum_exp(local_pes_30_22_io_out_sum_exp),
    .io_out_kv(local_pes_30_22_io_out_kv),
    .io_out_stage(local_pes_30_22_io_out_stage)
  );
  PE_1 local_pes_30_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_23_clock),
    .reset(local_pes_30_23_reset),
    .io_in_q(local_pes_30_23_io_in_q),
    .io_in_sum(local_pes_30_23_io_in_sum),
    .io_in_sum_exp(local_pes_30_23_io_in_sum_exp),
    .io_in_kv(local_pes_30_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_23_io_in_inv_sum),
    .io_in_stage(local_pes_30_23_io_in_stage),
    .io_out_q(local_pes_30_23_io_out_q),
    .io_out_sum(local_pes_30_23_io_out_sum),
    .io_out_sum_exp(local_pes_30_23_io_out_sum_exp),
    .io_out_kv(local_pes_30_23_io_out_kv),
    .io_out_stage(local_pes_30_23_io_out_stage)
  );
  PE_1 local_pes_30_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_24_clock),
    .reset(local_pes_30_24_reset),
    .io_in_q(local_pes_30_24_io_in_q),
    .io_in_sum(local_pes_30_24_io_in_sum),
    .io_in_sum_exp(local_pes_30_24_io_in_sum_exp),
    .io_in_kv(local_pes_30_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_24_io_in_inv_sum),
    .io_in_stage(local_pes_30_24_io_in_stage),
    .io_out_q(local_pes_30_24_io_out_q),
    .io_out_sum(local_pes_30_24_io_out_sum),
    .io_out_sum_exp(local_pes_30_24_io_out_sum_exp),
    .io_out_kv(local_pes_30_24_io_out_kv),
    .io_out_stage(local_pes_30_24_io_out_stage)
  );
  PE_1 local_pes_30_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_25_clock),
    .reset(local_pes_30_25_reset),
    .io_in_q(local_pes_30_25_io_in_q),
    .io_in_sum(local_pes_30_25_io_in_sum),
    .io_in_sum_exp(local_pes_30_25_io_in_sum_exp),
    .io_in_kv(local_pes_30_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_25_io_in_inv_sum),
    .io_in_stage(local_pes_30_25_io_in_stage),
    .io_out_q(local_pes_30_25_io_out_q),
    .io_out_sum(local_pes_30_25_io_out_sum),
    .io_out_sum_exp(local_pes_30_25_io_out_sum_exp),
    .io_out_kv(local_pes_30_25_io_out_kv),
    .io_out_stage(local_pes_30_25_io_out_stage)
  );
  PE_1 local_pes_30_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_26_clock),
    .reset(local_pes_30_26_reset),
    .io_in_q(local_pes_30_26_io_in_q),
    .io_in_sum(local_pes_30_26_io_in_sum),
    .io_in_sum_exp(local_pes_30_26_io_in_sum_exp),
    .io_in_kv(local_pes_30_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_26_io_in_inv_sum),
    .io_in_stage(local_pes_30_26_io_in_stage),
    .io_out_q(local_pes_30_26_io_out_q),
    .io_out_sum(local_pes_30_26_io_out_sum),
    .io_out_sum_exp(local_pes_30_26_io_out_sum_exp),
    .io_out_kv(local_pes_30_26_io_out_kv),
    .io_out_stage(local_pes_30_26_io_out_stage)
  );
  PE_1 local_pes_30_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_27_clock),
    .reset(local_pes_30_27_reset),
    .io_in_q(local_pes_30_27_io_in_q),
    .io_in_sum(local_pes_30_27_io_in_sum),
    .io_in_sum_exp(local_pes_30_27_io_in_sum_exp),
    .io_in_kv(local_pes_30_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_27_io_in_inv_sum),
    .io_in_stage(local_pes_30_27_io_in_stage),
    .io_out_q(local_pes_30_27_io_out_q),
    .io_out_sum(local_pes_30_27_io_out_sum),
    .io_out_sum_exp(local_pes_30_27_io_out_sum_exp),
    .io_out_kv(local_pes_30_27_io_out_kv),
    .io_out_stage(local_pes_30_27_io_out_stage)
  );
  PE_1 local_pes_30_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_28_clock),
    .reset(local_pes_30_28_reset),
    .io_in_q(local_pes_30_28_io_in_q),
    .io_in_sum(local_pes_30_28_io_in_sum),
    .io_in_sum_exp(local_pes_30_28_io_in_sum_exp),
    .io_in_kv(local_pes_30_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_28_io_in_inv_sum),
    .io_in_stage(local_pes_30_28_io_in_stage),
    .io_out_q(local_pes_30_28_io_out_q),
    .io_out_sum(local_pes_30_28_io_out_sum),
    .io_out_sum_exp(local_pes_30_28_io_out_sum_exp),
    .io_out_kv(local_pes_30_28_io_out_kv),
    .io_out_stage(local_pes_30_28_io_out_stage)
  );
  PE_1 local_pes_30_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_29_clock),
    .reset(local_pes_30_29_reset),
    .io_in_q(local_pes_30_29_io_in_q),
    .io_in_sum(local_pes_30_29_io_in_sum),
    .io_in_sum_exp(local_pes_30_29_io_in_sum_exp),
    .io_in_kv(local_pes_30_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_29_io_in_inv_sum),
    .io_in_stage(local_pes_30_29_io_in_stage),
    .io_out_q(local_pes_30_29_io_out_q),
    .io_out_sum(local_pes_30_29_io_out_sum),
    .io_out_sum_exp(local_pes_30_29_io_out_sum_exp),
    .io_out_kv(local_pes_30_29_io_out_kv),
    .io_out_stage(local_pes_30_29_io_out_stage)
  );
  PE_1 local_pes_30_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_30_clock),
    .reset(local_pes_30_30_reset),
    .io_in_q(local_pes_30_30_io_in_q),
    .io_in_sum(local_pes_30_30_io_in_sum),
    .io_in_sum_exp(local_pes_30_30_io_in_sum_exp),
    .io_in_kv(local_pes_30_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_30_io_in_inv_sum),
    .io_in_stage(local_pes_30_30_io_in_stage),
    .io_out_q(local_pes_30_30_io_out_q),
    .io_out_sum(local_pes_30_30_io_out_sum),
    .io_out_sum_exp(local_pes_30_30_io_out_sum_exp),
    .io_out_kv(local_pes_30_30_io_out_kv),
    .io_out_stage(local_pes_30_30_io_out_stage)
  );
  PE_1 local_pes_30_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_30_31_clock),
    .reset(local_pes_30_31_reset),
    .io_in_q(local_pes_30_31_io_in_q),
    .io_in_sum(local_pes_30_31_io_in_sum),
    .io_in_sum_exp(local_pes_30_31_io_in_sum_exp),
    .io_in_kv(local_pes_30_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_30_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_30_31_io_in_inv_sum),
    .io_in_stage(local_pes_30_31_io_in_stage),
    .io_out_q(local_pes_30_31_io_out_q),
    .io_out_sum(local_pes_30_31_io_out_sum),
    .io_out_sum_exp(local_pes_30_31_io_out_sum_exp),
    .io_out_kv(local_pes_30_31_io_out_kv),
    .io_out_stage(local_pes_30_31_io_out_stage)
  );
  PE local_pes_31_0 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_0_clock),
    .reset(local_pes_31_0_reset),
    .io_in_q(local_pes_31_0_io_in_q),
    .io_in_kv(local_pes_31_0_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_0_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_0_io_in_inv_sum),
    .io_in_stage(local_pes_31_0_io_in_stage),
    .io_out_q(local_pes_31_0_io_out_q),
    .io_out_sum(local_pes_31_0_io_out_sum),
    .io_out_kv(local_pes_31_0_io_out_kv),
    .io_out_stage(local_pes_31_0_io_out_stage)
  );
  PE_1 local_pes_31_1 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_1_clock),
    .reset(local_pes_31_1_reset),
    .io_in_q(local_pes_31_1_io_in_q),
    .io_in_sum(local_pes_31_1_io_in_sum),
    .io_in_sum_exp(local_pes_31_1_io_in_sum_exp),
    .io_in_kv(local_pes_31_1_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_1_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_1_io_in_inv_sum),
    .io_in_stage(local_pes_31_1_io_in_stage),
    .io_out_q(local_pes_31_1_io_out_q),
    .io_out_sum(local_pes_31_1_io_out_sum),
    .io_out_sum_exp(local_pes_31_1_io_out_sum_exp),
    .io_out_kv(local_pes_31_1_io_out_kv),
    .io_out_stage(local_pes_31_1_io_out_stage)
  );
  PE_1 local_pes_31_2 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_2_clock),
    .reset(local_pes_31_2_reset),
    .io_in_q(local_pes_31_2_io_in_q),
    .io_in_sum(local_pes_31_2_io_in_sum),
    .io_in_sum_exp(local_pes_31_2_io_in_sum_exp),
    .io_in_kv(local_pes_31_2_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_2_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_2_io_in_inv_sum),
    .io_in_stage(local_pes_31_2_io_in_stage),
    .io_out_q(local_pes_31_2_io_out_q),
    .io_out_sum(local_pes_31_2_io_out_sum),
    .io_out_sum_exp(local_pes_31_2_io_out_sum_exp),
    .io_out_kv(local_pes_31_2_io_out_kv),
    .io_out_stage(local_pes_31_2_io_out_stage)
  );
  PE_1 local_pes_31_3 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_3_clock),
    .reset(local_pes_31_3_reset),
    .io_in_q(local_pes_31_3_io_in_q),
    .io_in_sum(local_pes_31_3_io_in_sum),
    .io_in_sum_exp(local_pes_31_3_io_in_sum_exp),
    .io_in_kv(local_pes_31_3_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_3_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_3_io_in_inv_sum),
    .io_in_stage(local_pes_31_3_io_in_stage),
    .io_out_q(local_pes_31_3_io_out_q),
    .io_out_sum(local_pes_31_3_io_out_sum),
    .io_out_sum_exp(local_pes_31_3_io_out_sum_exp),
    .io_out_kv(local_pes_31_3_io_out_kv),
    .io_out_stage(local_pes_31_3_io_out_stage)
  );
  PE_1 local_pes_31_4 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_4_clock),
    .reset(local_pes_31_4_reset),
    .io_in_q(local_pes_31_4_io_in_q),
    .io_in_sum(local_pes_31_4_io_in_sum),
    .io_in_sum_exp(local_pes_31_4_io_in_sum_exp),
    .io_in_kv(local_pes_31_4_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_4_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_4_io_in_inv_sum),
    .io_in_stage(local_pes_31_4_io_in_stage),
    .io_out_q(local_pes_31_4_io_out_q),
    .io_out_sum(local_pes_31_4_io_out_sum),
    .io_out_sum_exp(local_pes_31_4_io_out_sum_exp),
    .io_out_kv(local_pes_31_4_io_out_kv),
    .io_out_stage(local_pes_31_4_io_out_stage)
  );
  PE_1 local_pes_31_5 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_5_clock),
    .reset(local_pes_31_5_reset),
    .io_in_q(local_pes_31_5_io_in_q),
    .io_in_sum(local_pes_31_5_io_in_sum),
    .io_in_sum_exp(local_pes_31_5_io_in_sum_exp),
    .io_in_kv(local_pes_31_5_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_5_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_5_io_in_inv_sum),
    .io_in_stage(local_pes_31_5_io_in_stage),
    .io_out_q(local_pes_31_5_io_out_q),
    .io_out_sum(local_pes_31_5_io_out_sum),
    .io_out_sum_exp(local_pes_31_5_io_out_sum_exp),
    .io_out_kv(local_pes_31_5_io_out_kv),
    .io_out_stage(local_pes_31_5_io_out_stage)
  );
  PE_1 local_pes_31_6 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_6_clock),
    .reset(local_pes_31_6_reset),
    .io_in_q(local_pes_31_6_io_in_q),
    .io_in_sum(local_pes_31_6_io_in_sum),
    .io_in_sum_exp(local_pes_31_6_io_in_sum_exp),
    .io_in_kv(local_pes_31_6_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_6_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_6_io_in_inv_sum),
    .io_in_stage(local_pes_31_6_io_in_stage),
    .io_out_q(local_pes_31_6_io_out_q),
    .io_out_sum(local_pes_31_6_io_out_sum),
    .io_out_sum_exp(local_pes_31_6_io_out_sum_exp),
    .io_out_kv(local_pes_31_6_io_out_kv),
    .io_out_stage(local_pes_31_6_io_out_stage)
  );
  PE_1 local_pes_31_7 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_7_clock),
    .reset(local_pes_31_7_reset),
    .io_in_q(local_pes_31_7_io_in_q),
    .io_in_sum(local_pes_31_7_io_in_sum),
    .io_in_sum_exp(local_pes_31_7_io_in_sum_exp),
    .io_in_kv(local_pes_31_7_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_7_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_7_io_in_inv_sum),
    .io_in_stage(local_pes_31_7_io_in_stage),
    .io_out_q(local_pes_31_7_io_out_q),
    .io_out_sum(local_pes_31_7_io_out_sum),
    .io_out_sum_exp(local_pes_31_7_io_out_sum_exp),
    .io_out_kv(local_pes_31_7_io_out_kv),
    .io_out_stage(local_pes_31_7_io_out_stage)
  );
  PE_1 local_pes_31_8 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_8_clock),
    .reset(local_pes_31_8_reset),
    .io_in_q(local_pes_31_8_io_in_q),
    .io_in_sum(local_pes_31_8_io_in_sum),
    .io_in_sum_exp(local_pes_31_8_io_in_sum_exp),
    .io_in_kv(local_pes_31_8_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_8_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_8_io_in_inv_sum),
    .io_in_stage(local_pes_31_8_io_in_stage),
    .io_out_q(local_pes_31_8_io_out_q),
    .io_out_sum(local_pes_31_8_io_out_sum),
    .io_out_sum_exp(local_pes_31_8_io_out_sum_exp),
    .io_out_kv(local_pes_31_8_io_out_kv),
    .io_out_stage(local_pes_31_8_io_out_stage)
  );
  PE_1 local_pes_31_9 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_9_clock),
    .reset(local_pes_31_9_reset),
    .io_in_q(local_pes_31_9_io_in_q),
    .io_in_sum(local_pes_31_9_io_in_sum),
    .io_in_sum_exp(local_pes_31_9_io_in_sum_exp),
    .io_in_kv(local_pes_31_9_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_9_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_9_io_in_inv_sum),
    .io_in_stage(local_pes_31_9_io_in_stage),
    .io_out_q(local_pes_31_9_io_out_q),
    .io_out_sum(local_pes_31_9_io_out_sum),
    .io_out_sum_exp(local_pes_31_9_io_out_sum_exp),
    .io_out_kv(local_pes_31_9_io_out_kv),
    .io_out_stage(local_pes_31_9_io_out_stage)
  );
  PE_1 local_pes_31_10 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_10_clock),
    .reset(local_pes_31_10_reset),
    .io_in_q(local_pes_31_10_io_in_q),
    .io_in_sum(local_pes_31_10_io_in_sum),
    .io_in_sum_exp(local_pes_31_10_io_in_sum_exp),
    .io_in_kv(local_pes_31_10_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_10_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_10_io_in_inv_sum),
    .io_in_stage(local_pes_31_10_io_in_stage),
    .io_out_q(local_pes_31_10_io_out_q),
    .io_out_sum(local_pes_31_10_io_out_sum),
    .io_out_sum_exp(local_pes_31_10_io_out_sum_exp),
    .io_out_kv(local_pes_31_10_io_out_kv),
    .io_out_stage(local_pes_31_10_io_out_stage)
  );
  PE_1 local_pes_31_11 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_11_clock),
    .reset(local_pes_31_11_reset),
    .io_in_q(local_pes_31_11_io_in_q),
    .io_in_sum(local_pes_31_11_io_in_sum),
    .io_in_sum_exp(local_pes_31_11_io_in_sum_exp),
    .io_in_kv(local_pes_31_11_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_11_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_11_io_in_inv_sum),
    .io_in_stage(local_pes_31_11_io_in_stage),
    .io_out_q(local_pes_31_11_io_out_q),
    .io_out_sum(local_pes_31_11_io_out_sum),
    .io_out_sum_exp(local_pes_31_11_io_out_sum_exp),
    .io_out_kv(local_pes_31_11_io_out_kv),
    .io_out_stage(local_pes_31_11_io_out_stage)
  );
  PE_1 local_pes_31_12 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_12_clock),
    .reset(local_pes_31_12_reset),
    .io_in_q(local_pes_31_12_io_in_q),
    .io_in_sum(local_pes_31_12_io_in_sum),
    .io_in_sum_exp(local_pes_31_12_io_in_sum_exp),
    .io_in_kv(local_pes_31_12_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_12_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_12_io_in_inv_sum),
    .io_in_stage(local_pes_31_12_io_in_stage),
    .io_out_q(local_pes_31_12_io_out_q),
    .io_out_sum(local_pes_31_12_io_out_sum),
    .io_out_sum_exp(local_pes_31_12_io_out_sum_exp),
    .io_out_kv(local_pes_31_12_io_out_kv),
    .io_out_stage(local_pes_31_12_io_out_stage)
  );
  PE_1 local_pes_31_13 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_13_clock),
    .reset(local_pes_31_13_reset),
    .io_in_q(local_pes_31_13_io_in_q),
    .io_in_sum(local_pes_31_13_io_in_sum),
    .io_in_sum_exp(local_pes_31_13_io_in_sum_exp),
    .io_in_kv(local_pes_31_13_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_13_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_13_io_in_inv_sum),
    .io_in_stage(local_pes_31_13_io_in_stage),
    .io_out_q(local_pes_31_13_io_out_q),
    .io_out_sum(local_pes_31_13_io_out_sum),
    .io_out_sum_exp(local_pes_31_13_io_out_sum_exp),
    .io_out_kv(local_pes_31_13_io_out_kv),
    .io_out_stage(local_pes_31_13_io_out_stage)
  );
  PE_1 local_pes_31_14 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_14_clock),
    .reset(local_pes_31_14_reset),
    .io_in_q(local_pes_31_14_io_in_q),
    .io_in_sum(local_pes_31_14_io_in_sum),
    .io_in_sum_exp(local_pes_31_14_io_in_sum_exp),
    .io_in_kv(local_pes_31_14_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_14_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_14_io_in_inv_sum),
    .io_in_stage(local_pes_31_14_io_in_stage),
    .io_out_q(local_pes_31_14_io_out_q),
    .io_out_sum(local_pes_31_14_io_out_sum),
    .io_out_sum_exp(local_pes_31_14_io_out_sum_exp),
    .io_out_kv(local_pes_31_14_io_out_kv),
    .io_out_stage(local_pes_31_14_io_out_stage)
  );
  PE_1 local_pes_31_15 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_15_clock),
    .reset(local_pes_31_15_reset),
    .io_in_q(local_pes_31_15_io_in_q),
    .io_in_sum(local_pes_31_15_io_in_sum),
    .io_in_sum_exp(local_pes_31_15_io_in_sum_exp),
    .io_in_kv(local_pes_31_15_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_15_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_15_io_in_inv_sum),
    .io_in_stage(local_pes_31_15_io_in_stage),
    .io_out_q(local_pes_31_15_io_out_q),
    .io_out_sum(local_pes_31_15_io_out_sum),
    .io_out_sum_exp(local_pes_31_15_io_out_sum_exp),
    .io_out_kv(local_pes_31_15_io_out_kv),
    .io_out_stage(local_pes_31_15_io_out_stage)
  );
  PE_1 local_pes_31_16 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_16_clock),
    .reset(local_pes_31_16_reset),
    .io_in_q(local_pes_31_16_io_in_q),
    .io_in_sum(local_pes_31_16_io_in_sum),
    .io_in_sum_exp(local_pes_31_16_io_in_sum_exp),
    .io_in_kv(local_pes_31_16_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_16_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_16_io_in_inv_sum),
    .io_in_stage(local_pes_31_16_io_in_stage),
    .io_out_q(local_pes_31_16_io_out_q),
    .io_out_sum(local_pes_31_16_io_out_sum),
    .io_out_sum_exp(local_pes_31_16_io_out_sum_exp),
    .io_out_kv(local_pes_31_16_io_out_kv),
    .io_out_stage(local_pes_31_16_io_out_stage)
  );
  PE_1 local_pes_31_17 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_17_clock),
    .reset(local_pes_31_17_reset),
    .io_in_q(local_pes_31_17_io_in_q),
    .io_in_sum(local_pes_31_17_io_in_sum),
    .io_in_sum_exp(local_pes_31_17_io_in_sum_exp),
    .io_in_kv(local_pes_31_17_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_17_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_17_io_in_inv_sum),
    .io_in_stage(local_pes_31_17_io_in_stage),
    .io_out_q(local_pes_31_17_io_out_q),
    .io_out_sum(local_pes_31_17_io_out_sum),
    .io_out_sum_exp(local_pes_31_17_io_out_sum_exp),
    .io_out_kv(local_pes_31_17_io_out_kv),
    .io_out_stage(local_pes_31_17_io_out_stage)
  );
  PE_1 local_pes_31_18 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_18_clock),
    .reset(local_pes_31_18_reset),
    .io_in_q(local_pes_31_18_io_in_q),
    .io_in_sum(local_pes_31_18_io_in_sum),
    .io_in_sum_exp(local_pes_31_18_io_in_sum_exp),
    .io_in_kv(local_pes_31_18_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_18_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_18_io_in_inv_sum),
    .io_in_stage(local_pes_31_18_io_in_stage),
    .io_out_q(local_pes_31_18_io_out_q),
    .io_out_sum(local_pes_31_18_io_out_sum),
    .io_out_sum_exp(local_pes_31_18_io_out_sum_exp),
    .io_out_kv(local_pes_31_18_io_out_kv),
    .io_out_stage(local_pes_31_18_io_out_stage)
  );
  PE_1 local_pes_31_19 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_19_clock),
    .reset(local_pes_31_19_reset),
    .io_in_q(local_pes_31_19_io_in_q),
    .io_in_sum(local_pes_31_19_io_in_sum),
    .io_in_sum_exp(local_pes_31_19_io_in_sum_exp),
    .io_in_kv(local_pes_31_19_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_19_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_19_io_in_inv_sum),
    .io_in_stage(local_pes_31_19_io_in_stage),
    .io_out_q(local_pes_31_19_io_out_q),
    .io_out_sum(local_pes_31_19_io_out_sum),
    .io_out_sum_exp(local_pes_31_19_io_out_sum_exp),
    .io_out_kv(local_pes_31_19_io_out_kv),
    .io_out_stage(local_pes_31_19_io_out_stage)
  );
  PE_1 local_pes_31_20 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_20_clock),
    .reset(local_pes_31_20_reset),
    .io_in_q(local_pes_31_20_io_in_q),
    .io_in_sum(local_pes_31_20_io_in_sum),
    .io_in_sum_exp(local_pes_31_20_io_in_sum_exp),
    .io_in_kv(local_pes_31_20_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_20_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_20_io_in_inv_sum),
    .io_in_stage(local_pes_31_20_io_in_stage),
    .io_out_q(local_pes_31_20_io_out_q),
    .io_out_sum(local_pes_31_20_io_out_sum),
    .io_out_sum_exp(local_pes_31_20_io_out_sum_exp),
    .io_out_kv(local_pes_31_20_io_out_kv),
    .io_out_stage(local_pes_31_20_io_out_stage)
  );
  PE_1 local_pes_31_21 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_21_clock),
    .reset(local_pes_31_21_reset),
    .io_in_q(local_pes_31_21_io_in_q),
    .io_in_sum(local_pes_31_21_io_in_sum),
    .io_in_sum_exp(local_pes_31_21_io_in_sum_exp),
    .io_in_kv(local_pes_31_21_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_21_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_21_io_in_inv_sum),
    .io_in_stage(local_pes_31_21_io_in_stage),
    .io_out_q(local_pes_31_21_io_out_q),
    .io_out_sum(local_pes_31_21_io_out_sum),
    .io_out_sum_exp(local_pes_31_21_io_out_sum_exp),
    .io_out_kv(local_pes_31_21_io_out_kv),
    .io_out_stage(local_pes_31_21_io_out_stage)
  );
  PE_1 local_pes_31_22 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_22_clock),
    .reset(local_pes_31_22_reset),
    .io_in_q(local_pes_31_22_io_in_q),
    .io_in_sum(local_pes_31_22_io_in_sum),
    .io_in_sum_exp(local_pes_31_22_io_in_sum_exp),
    .io_in_kv(local_pes_31_22_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_22_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_22_io_in_inv_sum),
    .io_in_stage(local_pes_31_22_io_in_stage),
    .io_out_q(local_pes_31_22_io_out_q),
    .io_out_sum(local_pes_31_22_io_out_sum),
    .io_out_sum_exp(local_pes_31_22_io_out_sum_exp),
    .io_out_kv(local_pes_31_22_io_out_kv),
    .io_out_stage(local_pes_31_22_io_out_stage)
  );
  PE_1 local_pes_31_23 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_23_clock),
    .reset(local_pes_31_23_reset),
    .io_in_q(local_pes_31_23_io_in_q),
    .io_in_sum(local_pes_31_23_io_in_sum),
    .io_in_sum_exp(local_pes_31_23_io_in_sum_exp),
    .io_in_kv(local_pes_31_23_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_23_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_23_io_in_inv_sum),
    .io_in_stage(local_pes_31_23_io_in_stage),
    .io_out_q(local_pes_31_23_io_out_q),
    .io_out_sum(local_pes_31_23_io_out_sum),
    .io_out_sum_exp(local_pes_31_23_io_out_sum_exp),
    .io_out_kv(local_pes_31_23_io_out_kv),
    .io_out_stage(local_pes_31_23_io_out_stage)
  );
  PE_1 local_pes_31_24 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_24_clock),
    .reset(local_pes_31_24_reset),
    .io_in_q(local_pes_31_24_io_in_q),
    .io_in_sum(local_pes_31_24_io_in_sum),
    .io_in_sum_exp(local_pes_31_24_io_in_sum_exp),
    .io_in_kv(local_pes_31_24_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_24_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_24_io_in_inv_sum),
    .io_in_stage(local_pes_31_24_io_in_stage),
    .io_out_q(local_pes_31_24_io_out_q),
    .io_out_sum(local_pes_31_24_io_out_sum),
    .io_out_sum_exp(local_pes_31_24_io_out_sum_exp),
    .io_out_kv(local_pes_31_24_io_out_kv),
    .io_out_stage(local_pes_31_24_io_out_stage)
  );
  PE_1 local_pes_31_25 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_25_clock),
    .reset(local_pes_31_25_reset),
    .io_in_q(local_pes_31_25_io_in_q),
    .io_in_sum(local_pes_31_25_io_in_sum),
    .io_in_sum_exp(local_pes_31_25_io_in_sum_exp),
    .io_in_kv(local_pes_31_25_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_25_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_25_io_in_inv_sum),
    .io_in_stage(local_pes_31_25_io_in_stage),
    .io_out_q(local_pes_31_25_io_out_q),
    .io_out_sum(local_pes_31_25_io_out_sum),
    .io_out_sum_exp(local_pes_31_25_io_out_sum_exp),
    .io_out_kv(local_pes_31_25_io_out_kv),
    .io_out_stage(local_pes_31_25_io_out_stage)
  );
  PE_1 local_pes_31_26 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_26_clock),
    .reset(local_pes_31_26_reset),
    .io_in_q(local_pes_31_26_io_in_q),
    .io_in_sum(local_pes_31_26_io_in_sum),
    .io_in_sum_exp(local_pes_31_26_io_in_sum_exp),
    .io_in_kv(local_pes_31_26_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_26_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_26_io_in_inv_sum),
    .io_in_stage(local_pes_31_26_io_in_stage),
    .io_out_q(local_pes_31_26_io_out_q),
    .io_out_sum(local_pes_31_26_io_out_sum),
    .io_out_sum_exp(local_pes_31_26_io_out_sum_exp),
    .io_out_kv(local_pes_31_26_io_out_kv),
    .io_out_stage(local_pes_31_26_io_out_stage)
  );
  PE_1 local_pes_31_27 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_27_clock),
    .reset(local_pes_31_27_reset),
    .io_in_q(local_pes_31_27_io_in_q),
    .io_in_sum(local_pes_31_27_io_in_sum),
    .io_in_sum_exp(local_pes_31_27_io_in_sum_exp),
    .io_in_kv(local_pes_31_27_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_27_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_27_io_in_inv_sum),
    .io_in_stage(local_pes_31_27_io_in_stage),
    .io_out_q(local_pes_31_27_io_out_q),
    .io_out_sum(local_pes_31_27_io_out_sum),
    .io_out_sum_exp(local_pes_31_27_io_out_sum_exp),
    .io_out_kv(local_pes_31_27_io_out_kv),
    .io_out_stage(local_pes_31_27_io_out_stage)
  );
  PE_1 local_pes_31_28 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_28_clock),
    .reset(local_pes_31_28_reset),
    .io_in_q(local_pes_31_28_io_in_q),
    .io_in_sum(local_pes_31_28_io_in_sum),
    .io_in_sum_exp(local_pes_31_28_io_in_sum_exp),
    .io_in_kv(local_pes_31_28_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_28_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_28_io_in_inv_sum),
    .io_in_stage(local_pes_31_28_io_in_stage),
    .io_out_q(local_pes_31_28_io_out_q),
    .io_out_sum(local_pes_31_28_io_out_sum),
    .io_out_sum_exp(local_pes_31_28_io_out_sum_exp),
    .io_out_kv(local_pes_31_28_io_out_kv),
    .io_out_stage(local_pes_31_28_io_out_stage)
  );
  PE_1 local_pes_31_29 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_29_clock),
    .reset(local_pes_31_29_reset),
    .io_in_q(local_pes_31_29_io_in_q),
    .io_in_sum(local_pes_31_29_io_in_sum),
    .io_in_sum_exp(local_pes_31_29_io_in_sum_exp),
    .io_in_kv(local_pes_31_29_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_29_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_29_io_in_inv_sum),
    .io_in_stage(local_pes_31_29_io_in_stage),
    .io_out_q(local_pes_31_29_io_out_q),
    .io_out_sum(local_pes_31_29_io_out_sum),
    .io_out_sum_exp(local_pes_31_29_io_out_sum_exp),
    .io_out_kv(local_pes_31_29_io_out_kv),
    .io_out_stage(local_pes_31_29_io_out_stage)
  );
  PE_1 local_pes_31_30 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_30_clock),
    .reset(local_pes_31_30_reset),
    .io_in_q(local_pes_31_30_io_in_q),
    .io_in_sum(local_pes_31_30_io_in_sum),
    .io_in_sum_exp(local_pes_31_30_io_in_sum_exp),
    .io_in_kv(local_pes_31_30_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_30_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_30_io_in_inv_sum),
    .io_in_stage(local_pes_31_30_io_in_stage),
    .io_out_q(local_pes_31_30_io_out_q),
    .io_out_sum(local_pes_31_30_io_out_sum),
    .io_out_sum_exp(local_pes_31_30_io_out_sum_exp),
    .io_out_kv(local_pes_31_30_io_out_kv),
    .io_out_stage(local_pes_31_30_io_out_stage)
  );
  PE_1 local_pes_31_31 ( // @[PEArray.scala 23:49]
    .clock(local_pes_31_31_clock),
    .reset(local_pes_31_31_reset),
    .io_in_q(local_pes_31_31_io_in_q),
    .io_in_sum(local_pes_31_31_io_in_sum),
    .io_in_sum_exp(local_pes_31_31_io_in_sum_exp),
    .io_in_kv(local_pes_31_31_io_in_kv),
    .io_in_inv_sum_exp(local_pes_31_31_io_in_inv_sum_exp),
    .io_in_inv_sum(local_pes_31_31_io_in_inv_sum),
    .io_in_stage(local_pes_31_31_io_in_stage),
    .io_out_q(local_pes_31_31_io_out_q),
    .io_out_sum(local_pes_31_31_io_out_sum),
    .io_out_sum_exp(local_pes_31_31_io_out_sum_exp),
    .io_out_kv(local_pes_31_31_io_out_kv),
    .io_out_stage(local_pes_31_31_io_out_stage)
  );
  PE_1 global_col_pes_0_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_0_0_clock),
    .reset(global_col_pes_0_0_reset),
    .io_in_q(global_col_pes_0_0_io_in_q),
    .io_in_sum(global_col_pes_0_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_0_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_0_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_0_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_0_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_0_0_io_in_stage),
    .io_out_q(global_col_pes_0_0_io_out_q),
    .io_out_sum(global_col_pes_0_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_0_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_0_0_io_out_kv),
    .io_out_stage(global_col_pes_0_0_io_out_stage)
  );
  PE_1 global_col_pes_1_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_1_0_clock),
    .reset(global_col_pes_1_0_reset),
    .io_in_q(global_col_pes_1_0_io_in_q),
    .io_in_sum(global_col_pes_1_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_1_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_1_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_1_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_1_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_1_0_io_in_stage),
    .io_out_q(global_col_pes_1_0_io_out_q),
    .io_out_sum(global_col_pes_1_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_1_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_1_0_io_out_kv),
    .io_out_stage(global_col_pes_1_0_io_out_stage)
  );
  PE_1 global_col_pes_2_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_2_0_clock),
    .reset(global_col_pes_2_0_reset),
    .io_in_q(global_col_pes_2_0_io_in_q),
    .io_in_sum(global_col_pes_2_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_2_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_2_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_2_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_2_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_2_0_io_in_stage),
    .io_out_q(global_col_pes_2_0_io_out_q),
    .io_out_sum(global_col_pes_2_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_2_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_2_0_io_out_kv),
    .io_out_stage(global_col_pes_2_0_io_out_stage)
  );
  PE_1 global_col_pes_3_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_3_0_clock),
    .reset(global_col_pes_3_0_reset),
    .io_in_q(global_col_pes_3_0_io_in_q),
    .io_in_sum(global_col_pes_3_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_3_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_3_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_3_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_3_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_3_0_io_in_stage),
    .io_out_q(global_col_pes_3_0_io_out_q),
    .io_out_sum(global_col_pes_3_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_3_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_3_0_io_out_kv),
    .io_out_stage(global_col_pes_3_0_io_out_stage)
  );
  PE_1 global_col_pes_4_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_4_0_clock),
    .reset(global_col_pes_4_0_reset),
    .io_in_q(global_col_pes_4_0_io_in_q),
    .io_in_sum(global_col_pes_4_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_4_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_4_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_4_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_4_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_4_0_io_in_stage),
    .io_out_q(global_col_pes_4_0_io_out_q),
    .io_out_sum(global_col_pes_4_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_4_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_4_0_io_out_kv),
    .io_out_stage(global_col_pes_4_0_io_out_stage)
  );
  PE_1 global_col_pes_5_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_5_0_clock),
    .reset(global_col_pes_5_0_reset),
    .io_in_q(global_col_pes_5_0_io_in_q),
    .io_in_sum(global_col_pes_5_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_5_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_5_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_5_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_5_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_5_0_io_in_stage),
    .io_out_q(global_col_pes_5_0_io_out_q),
    .io_out_sum(global_col_pes_5_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_5_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_5_0_io_out_kv),
    .io_out_stage(global_col_pes_5_0_io_out_stage)
  );
  PE_1 global_col_pes_6_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_6_0_clock),
    .reset(global_col_pes_6_0_reset),
    .io_in_q(global_col_pes_6_0_io_in_q),
    .io_in_sum(global_col_pes_6_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_6_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_6_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_6_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_6_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_6_0_io_in_stage),
    .io_out_q(global_col_pes_6_0_io_out_q),
    .io_out_sum(global_col_pes_6_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_6_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_6_0_io_out_kv),
    .io_out_stage(global_col_pes_6_0_io_out_stage)
  );
  PE_1 global_col_pes_7_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_7_0_clock),
    .reset(global_col_pes_7_0_reset),
    .io_in_q(global_col_pes_7_0_io_in_q),
    .io_in_sum(global_col_pes_7_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_7_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_7_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_7_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_7_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_7_0_io_in_stage),
    .io_out_q(global_col_pes_7_0_io_out_q),
    .io_out_sum(global_col_pes_7_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_7_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_7_0_io_out_kv),
    .io_out_stage(global_col_pes_7_0_io_out_stage)
  );
  PE_1 global_col_pes_8_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_8_0_clock),
    .reset(global_col_pes_8_0_reset),
    .io_in_q(global_col_pes_8_0_io_in_q),
    .io_in_sum(global_col_pes_8_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_8_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_8_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_8_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_8_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_8_0_io_in_stage),
    .io_out_q(global_col_pes_8_0_io_out_q),
    .io_out_sum(global_col_pes_8_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_8_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_8_0_io_out_kv),
    .io_out_stage(global_col_pes_8_0_io_out_stage)
  );
  PE_1 global_col_pes_9_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_9_0_clock),
    .reset(global_col_pes_9_0_reset),
    .io_in_q(global_col_pes_9_0_io_in_q),
    .io_in_sum(global_col_pes_9_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_9_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_9_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_9_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_9_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_9_0_io_in_stage),
    .io_out_q(global_col_pes_9_0_io_out_q),
    .io_out_sum(global_col_pes_9_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_9_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_9_0_io_out_kv),
    .io_out_stage(global_col_pes_9_0_io_out_stage)
  );
  PE_1 global_col_pes_10_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_10_0_clock),
    .reset(global_col_pes_10_0_reset),
    .io_in_q(global_col_pes_10_0_io_in_q),
    .io_in_sum(global_col_pes_10_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_10_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_10_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_10_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_10_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_10_0_io_in_stage),
    .io_out_q(global_col_pes_10_0_io_out_q),
    .io_out_sum(global_col_pes_10_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_10_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_10_0_io_out_kv),
    .io_out_stage(global_col_pes_10_0_io_out_stage)
  );
  PE_1 global_col_pes_11_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_11_0_clock),
    .reset(global_col_pes_11_0_reset),
    .io_in_q(global_col_pes_11_0_io_in_q),
    .io_in_sum(global_col_pes_11_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_11_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_11_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_11_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_11_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_11_0_io_in_stage),
    .io_out_q(global_col_pes_11_0_io_out_q),
    .io_out_sum(global_col_pes_11_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_11_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_11_0_io_out_kv),
    .io_out_stage(global_col_pes_11_0_io_out_stage)
  );
  PE_1 global_col_pes_12_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_12_0_clock),
    .reset(global_col_pes_12_0_reset),
    .io_in_q(global_col_pes_12_0_io_in_q),
    .io_in_sum(global_col_pes_12_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_12_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_12_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_12_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_12_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_12_0_io_in_stage),
    .io_out_q(global_col_pes_12_0_io_out_q),
    .io_out_sum(global_col_pes_12_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_12_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_12_0_io_out_kv),
    .io_out_stage(global_col_pes_12_0_io_out_stage)
  );
  PE_1 global_col_pes_13_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_13_0_clock),
    .reset(global_col_pes_13_0_reset),
    .io_in_q(global_col_pes_13_0_io_in_q),
    .io_in_sum(global_col_pes_13_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_13_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_13_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_13_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_13_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_13_0_io_in_stage),
    .io_out_q(global_col_pes_13_0_io_out_q),
    .io_out_sum(global_col_pes_13_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_13_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_13_0_io_out_kv),
    .io_out_stage(global_col_pes_13_0_io_out_stage)
  );
  PE_1 global_col_pes_14_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_14_0_clock),
    .reset(global_col_pes_14_0_reset),
    .io_in_q(global_col_pes_14_0_io_in_q),
    .io_in_sum(global_col_pes_14_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_14_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_14_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_14_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_14_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_14_0_io_in_stage),
    .io_out_q(global_col_pes_14_0_io_out_q),
    .io_out_sum(global_col_pes_14_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_14_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_14_0_io_out_kv),
    .io_out_stage(global_col_pes_14_0_io_out_stage)
  );
  PE_1 global_col_pes_15_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_15_0_clock),
    .reset(global_col_pes_15_0_reset),
    .io_in_q(global_col_pes_15_0_io_in_q),
    .io_in_sum(global_col_pes_15_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_15_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_15_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_15_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_15_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_15_0_io_in_stage),
    .io_out_q(global_col_pes_15_0_io_out_q),
    .io_out_sum(global_col_pes_15_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_15_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_15_0_io_out_kv),
    .io_out_stage(global_col_pes_15_0_io_out_stage)
  );
  PE_1 global_col_pes_16_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_16_0_clock),
    .reset(global_col_pes_16_0_reset),
    .io_in_q(global_col_pes_16_0_io_in_q),
    .io_in_sum(global_col_pes_16_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_16_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_16_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_16_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_16_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_16_0_io_in_stage),
    .io_out_q(global_col_pes_16_0_io_out_q),
    .io_out_sum(global_col_pes_16_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_16_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_16_0_io_out_kv),
    .io_out_stage(global_col_pes_16_0_io_out_stage)
  );
  PE_1 global_col_pes_17_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_17_0_clock),
    .reset(global_col_pes_17_0_reset),
    .io_in_q(global_col_pes_17_0_io_in_q),
    .io_in_sum(global_col_pes_17_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_17_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_17_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_17_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_17_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_17_0_io_in_stage),
    .io_out_q(global_col_pes_17_0_io_out_q),
    .io_out_sum(global_col_pes_17_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_17_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_17_0_io_out_kv),
    .io_out_stage(global_col_pes_17_0_io_out_stage)
  );
  PE_1 global_col_pes_18_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_18_0_clock),
    .reset(global_col_pes_18_0_reset),
    .io_in_q(global_col_pes_18_0_io_in_q),
    .io_in_sum(global_col_pes_18_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_18_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_18_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_18_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_18_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_18_0_io_in_stage),
    .io_out_q(global_col_pes_18_0_io_out_q),
    .io_out_sum(global_col_pes_18_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_18_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_18_0_io_out_kv),
    .io_out_stage(global_col_pes_18_0_io_out_stage)
  );
  PE_1 global_col_pes_19_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_19_0_clock),
    .reset(global_col_pes_19_0_reset),
    .io_in_q(global_col_pes_19_0_io_in_q),
    .io_in_sum(global_col_pes_19_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_19_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_19_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_19_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_19_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_19_0_io_in_stage),
    .io_out_q(global_col_pes_19_0_io_out_q),
    .io_out_sum(global_col_pes_19_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_19_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_19_0_io_out_kv),
    .io_out_stage(global_col_pes_19_0_io_out_stage)
  );
  PE_1 global_col_pes_20_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_20_0_clock),
    .reset(global_col_pes_20_0_reset),
    .io_in_q(global_col_pes_20_0_io_in_q),
    .io_in_sum(global_col_pes_20_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_20_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_20_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_20_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_20_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_20_0_io_in_stage),
    .io_out_q(global_col_pes_20_0_io_out_q),
    .io_out_sum(global_col_pes_20_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_20_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_20_0_io_out_kv),
    .io_out_stage(global_col_pes_20_0_io_out_stage)
  );
  PE_1 global_col_pes_21_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_21_0_clock),
    .reset(global_col_pes_21_0_reset),
    .io_in_q(global_col_pes_21_0_io_in_q),
    .io_in_sum(global_col_pes_21_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_21_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_21_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_21_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_21_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_21_0_io_in_stage),
    .io_out_q(global_col_pes_21_0_io_out_q),
    .io_out_sum(global_col_pes_21_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_21_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_21_0_io_out_kv),
    .io_out_stage(global_col_pes_21_0_io_out_stage)
  );
  PE_1 global_col_pes_22_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_22_0_clock),
    .reset(global_col_pes_22_0_reset),
    .io_in_q(global_col_pes_22_0_io_in_q),
    .io_in_sum(global_col_pes_22_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_22_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_22_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_22_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_22_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_22_0_io_in_stage),
    .io_out_q(global_col_pes_22_0_io_out_q),
    .io_out_sum(global_col_pes_22_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_22_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_22_0_io_out_kv),
    .io_out_stage(global_col_pes_22_0_io_out_stage)
  );
  PE_1 global_col_pes_23_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_23_0_clock),
    .reset(global_col_pes_23_0_reset),
    .io_in_q(global_col_pes_23_0_io_in_q),
    .io_in_sum(global_col_pes_23_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_23_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_23_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_23_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_23_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_23_0_io_in_stage),
    .io_out_q(global_col_pes_23_0_io_out_q),
    .io_out_sum(global_col_pes_23_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_23_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_23_0_io_out_kv),
    .io_out_stage(global_col_pes_23_0_io_out_stage)
  );
  PE_1 global_col_pes_24_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_24_0_clock),
    .reset(global_col_pes_24_0_reset),
    .io_in_q(global_col_pes_24_0_io_in_q),
    .io_in_sum(global_col_pes_24_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_24_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_24_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_24_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_24_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_24_0_io_in_stage),
    .io_out_q(global_col_pes_24_0_io_out_q),
    .io_out_sum(global_col_pes_24_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_24_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_24_0_io_out_kv),
    .io_out_stage(global_col_pes_24_0_io_out_stage)
  );
  PE_1 global_col_pes_25_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_25_0_clock),
    .reset(global_col_pes_25_0_reset),
    .io_in_q(global_col_pes_25_0_io_in_q),
    .io_in_sum(global_col_pes_25_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_25_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_25_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_25_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_25_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_25_0_io_in_stage),
    .io_out_q(global_col_pes_25_0_io_out_q),
    .io_out_sum(global_col_pes_25_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_25_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_25_0_io_out_kv),
    .io_out_stage(global_col_pes_25_0_io_out_stage)
  );
  PE_1 global_col_pes_26_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_26_0_clock),
    .reset(global_col_pes_26_0_reset),
    .io_in_q(global_col_pes_26_0_io_in_q),
    .io_in_sum(global_col_pes_26_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_26_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_26_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_26_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_26_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_26_0_io_in_stage),
    .io_out_q(global_col_pes_26_0_io_out_q),
    .io_out_sum(global_col_pes_26_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_26_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_26_0_io_out_kv),
    .io_out_stage(global_col_pes_26_0_io_out_stage)
  );
  PE_1 global_col_pes_27_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_27_0_clock),
    .reset(global_col_pes_27_0_reset),
    .io_in_q(global_col_pes_27_0_io_in_q),
    .io_in_sum(global_col_pes_27_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_27_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_27_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_27_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_27_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_27_0_io_in_stage),
    .io_out_q(global_col_pes_27_0_io_out_q),
    .io_out_sum(global_col_pes_27_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_27_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_27_0_io_out_kv),
    .io_out_stage(global_col_pes_27_0_io_out_stage)
  );
  PE_1 global_col_pes_28_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_28_0_clock),
    .reset(global_col_pes_28_0_reset),
    .io_in_q(global_col_pes_28_0_io_in_q),
    .io_in_sum(global_col_pes_28_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_28_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_28_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_28_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_28_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_28_0_io_in_stage),
    .io_out_q(global_col_pes_28_0_io_out_q),
    .io_out_sum(global_col_pes_28_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_28_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_28_0_io_out_kv),
    .io_out_stage(global_col_pes_28_0_io_out_stage)
  );
  PE_1 global_col_pes_29_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_29_0_clock),
    .reset(global_col_pes_29_0_reset),
    .io_in_q(global_col_pes_29_0_io_in_q),
    .io_in_sum(global_col_pes_29_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_29_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_29_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_29_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_29_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_29_0_io_in_stage),
    .io_out_q(global_col_pes_29_0_io_out_q),
    .io_out_sum(global_col_pes_29_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_29_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_29_0_io_out_kv),
    .io_out_stage(global_col_pes_29_0_io_out_stage)
  );
  PE_1 global_col_pes_30_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_30_0_clock),
    .reset(global_col_pes_30_0_reset),
    .io_in_q(global_col_pes_30_0_io_in_q),
    .io_in_sum(global_col_pes_30_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_30_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_30_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_30_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_30_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_30_0_io_in_stage),
    .io_out_q(global_col_pes_30_0_io_out_q),
    .io_out_sum(global_col_pes_30_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_30_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_30_0_io_out_kv),
    .io_out_stage(global_col_pes_30_0_io_out_stage)
  );
  PE_1 global_col_pes_31_0 ( // @[PEArray.scala 26:50]
    .clock(global_col_pes_31_0_clock),
    .reset(global_col_pes_31_0_reset),
    .io_in_q(global_col_pes_31_0_io_in_q),
    .io_in_sum(global_col_pes_31_0_io_in_sum),
    .io_in_sum_exp(global_col_pes_31_0_io_in_sum_exp),
    .io_in_kv(global_col_pes_31_0_io_in_kv),
    .io_in_inv_sum_exp(global_col_pes_31_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_col_pes_31_0_io_in_inv_sum),
    .io_in_stage(global_col_pes_31_0_io_in_stage),
    .io_out_q(global_col_pes_31_0_io_out_q),
    .io_out_sum(global_col_pes_31_0_io_out_sum),
    .io_out_sum_exp(global_col_pes_31_0_io_out_sum_exp),
    .io_out_kv(global_col_pes_31_0_io_out_kv),
    .io_out_stage(global_col_pes_31_0_io_out_stage)
  );
  PE global_row_pes_0_0 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_0_clock),
    .reset(global_row_pes_0_0_reset),
    .io_in_q(global_row_pes_0_0_io_in_q),
    .io_in_kv(global_row_pes_0_0_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_0_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_0_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_0_io_in_stage),
    .io_out_q(global_row_pes_0_0_io_out_q),
    .io_out_sum(global_row_pes_0_0_io_out_sum),
    .io_out_kv(global_row_pes_0_0_io_out_kv),
    .io_out_stage(global_row_pes_0_0_io_out_stage)
  );
  PE_1 global_row_pes_0_1 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_1_clock),
    .reset(global_row_pes_0_1_reset),
    .io_in_q(global_row_pes_0_1_io_in_q),
    .io_in_sum(global_row_pes_0_1_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_1_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_1_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_1_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_1_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_1_io_in_stage),
    .io_out_q(global_row_pes_0_1_io_out_q),
    .io_out_sum(global_row_pes_0_1_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_1_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_1_io_out_kv),
    .io_out_stage(global_row_pes_0_1_io_out_stage)
  );
  PE_1 global_row_pes_0_2 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_2_clock),
    .reset(global_row_pes_0_2_reset),
    .io_in_q(global_row_pes_0_2_io_in_q),
    .io_in_sum(global_row_pes_0_2_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_2_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_2_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_2_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_2_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_2_io_in_stage),
    .io_out_q(global_row_pes_0_2_io_out_q),
    .io_out_sum(global_row_pes_0_2_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_2_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_2_io_out_kv),
    .io_out_stage(global_row_pes_0_2_io_out_stage)
  );
  PE_1 global_row_pes_0_3 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_3_clock),
    .reset(global_row_pes_0_3_reset),
    .io_in_q(global_row_pes_0_3_io_in_q),
    .io_in_sum(global_row_pes_0_3_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_3_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_3_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_3_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_3_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_3_io_in_stage),
    .io_out_q(global_row_pes_0_3_io_out_q),
    .io_out_sum(global_row_pes_0_3_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_3_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_3_io_out_kv),
    .io_out_stage(global_row_pes_0_3_io_out_stage)
  );
  PE_1 global_row_pes_0_4 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_4_clock),
    .reset(global_row_pes_0_4_reset),
    .io_in_q(global_row_pes_0_4_io_in_q),
    .io_in_sum(global_row_pes_0_4_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_4_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_4_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_4_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_4_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_4_io_in_stage),
    .io_out_q(global_row_pes_0_4_io_out_q),
    .io_out_sum(global_row_pes_0_4_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_4_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_4_io_out_kv),
    .io_out_stage(global_row_pes_0_4_io_out_stage)
  );
  PE_1 global_row_pes_0_5 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_5_clock),
    .reset(global_row_pes_0_5_reset),
    .io_in_q(global_row_pes_0_5_io_in_q),
    .io_in_sum(global_row_pes_0_5_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_5_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_5_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_5_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_5_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_5_io_in_stage),
    .io_out_q(global_row_pes_0_5_io_out_q),
    .io_out_sum(global_row_pes_0_5_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_5_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_5_io_out_kv),
    .io_out_stage(global_row_pes_0_5_io_out_stage)
  );
  PE_1 global_row_pes_0_6 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_6_clock),
    .reset(global_row_pes_0_6_reset),
    .io_in_q(global_row_pes_0_6_io_in_q),
    .io_in_sum(global_row_pes_0_6_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_6_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_6_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_6_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_6_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_6_io_in_stage),
    .io_out_q(global_row_pes_0_6_io_out_q),
    .io_out_sum(global_row_pes_0_6_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_6_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_6_io_out_kv),
    .io_out_stage(global_row_pes_0_6_io_out_stage)
  );
  PE_1 global_row_pes_0_7 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_7_clock),
    .reset(global_row_pes_0_7_reset),
    .io_in_q(global_row_pes_0_7_io_in_q),
    .io_in_sum(global_row_pes_0_7_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_7_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_7_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_7_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_7_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_7_io_in_stage),
    .io_out_q(global_row_pes_0_7_io_out_q),
    .io_out_sum(global_row_pes_0_7_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_7_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_7_io_out_kv),
    .io_out_stage(global_row_pes_0_7_io_out_stage)
  );
  PE_1 global_row_pes_0_8 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_8_clock),
    .reset(global_row_pes_0_8_reset),
    .io_in_q(global_row_pes_0_8_io_in_q),
    .io_in_sum(global_row_pes_0_8_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_8_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_8_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_8_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_8_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_8_io_in_stage),
    .io_out_q(global_row_pes_0_8_io_out_q),
    .io_out_sum(global_row_pes_0_8_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_8_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_8_io_out_kv),
    .io_out_stage(global_row_pes_0_8_io_out_stage)
  );
  PE_1 global_row_pes_0_9 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_9_clock),
    .reset(global_row_pes_0_9_reset),
    .io_in_q(global_row_pes_0_9_io_in_q),
    .io_in_sum(global_row_pes_0_9_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_9_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_9_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_9_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_9_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_9_io_in_stage),
    .io_out_q(global_row_pes_0_9_io_out_q),
    .io_out_sum(global_row_pes_0_9_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_9_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_9_io_out_kv),
    .io_out_stage(global_row_pes_0_9_io_out_stage)
  );
  PE_1 global_row_pes_0_10 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_10_clock),
    .reset(global_row_pes_0_10_reset),
    .io_in_q(global_row_pes_0_10_io_in_q),
    .io_in_sum(global_row_pes_0_10_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_10_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_10_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_10_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_10_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_10_io_in_stage),
    .io_out_q(global_row_pes_0_10_io_out_q),
    .io_out_sum(global_row_pes_0_10_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_10_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_10_io_out_kv),
    .io_out_stage(global_row_pes_0_10_io_out_stage)
  );
  PE_1 global_row_pes_0_11 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_11_clock),
    .reset(global_row_pes_0_11_reset),
    .io_in_q(global_row_pes_0_11_io_in_q),
    .io_in_sum(global_row_pes_0_11_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_11_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_11_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_11_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_11_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_11_io_in_stage),
    .io_out_q(global_row_pes_0_11_io_out_q),
    .io_out_sum(global_row_pes_0_11_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_11_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_11_io_out_kv),
    .io_out_stage(global_row_pes_0_11_io_out_stage)
  );
  PE_1 global_row_pes_0_12 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_12_clock),
    .reset(global_row_pes_0_12_reset),
    .io_in_q(global_row_pes_0_12_io_in_q),
    .io_in_sum(global_row_pes_0_12_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_12_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_12_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_12_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_12_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_12_io_in_stage),
    .io_out_q(global_row_pes_0_12_io_out_q),
    .io_out_sum(global_row_pes_0_12_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_12_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_12_io_out_kv),
    .io_out_stage(global_row_pes_0_12_io_out_stage)
  );
  PE_1 global_row_pes_0_13 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_13_clock),
    .reset(global_row_pes_0_13_reset),
    .io_in_q(global_row_pes_0_13_io_in_q),
    .io_in_sum(global_row_pes_0_13_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_13_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_13_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_13_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_13_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_13_io_in_stage),
    .io_out_q(global_row_pes_0_13_io_out_q),
    .io_out_sum(global_row_pes_0_13_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_13_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_13_io_out_kv),
    .io_out_stage(global_row_pes_0_13_io_out_stage)
  );
  PE_1 global_row_pes_0_14 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_14_clock),
    .reset(global_row_pes_0_14_reset),
    .io_in_q(global_row_pes_0_14_io_in_q),
    .io_in_sum(global_row_pes_0_14_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_14_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_14_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_14_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_14_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_14_io_in_stage),
    .io_out_q(global_row_pes_0_14_io_out_q),
    .io_out_sum(global_row_pes_0_14_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_14_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_14_io_out_kv),
    .io_out_stage(global_row_pes_0_14_io_out_stage)
  );
  PE_1 global_row_pes_0_15 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_15_clock),
    .reset(global_row_pes_0_15_reset),
    .io_in_q(global_row_pes_0_15_io_in_q),
    .io_in_sum(global_row_pes_0_15_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_15_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_15_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_15_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_15_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_15_io_in_stage),
    .io_out_q(global_row_pes_0_15_io_out_q),
    .io_out_sum(global_row_pes_0_15_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_15_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_15_io_out_kv),
    .io_out_stage(global_row_pes_0_15_io_out_stage)
  );
  PE_1 global_row_pes_0_16 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_16_clock),
    .reset(global_row_pes_0_16_reset),
    .io_in_q(global_row_pes_0_16_io_in_q),
    .io_in_sum(global_row_pes_0_16_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_16_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_16_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_16_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_16_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_16_io_in_stage),
    .io_out_q(global_row_pes_0_16_io_out_q),
    .io_out_sum(global_row_pes_0_16_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_16_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_16_io_out_kv),
    .io_out_stage(global_row_pes_0_16_io_out_stage)
  );
  PE_1 global_row_pes_0_17 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_17_clock),
    .reset(global_row_pes_0_17_reset),
    .io_in_q(global_row_pes_0_17_io_in_q),
    .io_in_sum(global_row_pes_0_17_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_17_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_17_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_17_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_17_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_17_io_in_stage),
    .io_out_q(global_row_pes_0_17_io_out_q),
    .io_out_sum(global_row_pes_0_17_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_17_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_17_io_out_kv),
    .io_out_stage(global_row_pes_0_17_io_out_stage)
  );
  PE_1 global_row_pes_0_18 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_18_clock),
    .reset(global_row_pes_0_18_reset),
    .io_in_q(global_row_pes_0_18_io_in_q),
    .io_in_sum(global_row_pes_0_18_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_18_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_18_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_18_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_18_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_18_io_in_stage),
    .io_out_q(global_row_pes_0_18_io_out_q),
    .io_out_sum(global_row_pes_0_18_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_18_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_18_io_out_kv),
    .io_out_stage(global_row_pes_0_18_io_out_stage)
  );
  PE_1 global_row_pes_0_19 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_19_clock),
    .reset(global_row_pes_0_19_reset),
    .io_in_q(global_row_pes_0_19_io_in_q),
    .io_in_sum(global_row_pes_0_19_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_19_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_19_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_19_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_19_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_19_io_in_stage),
    .io_out_q(global_row_pes_0_19_io_out_q),
    .io_out_sum(global_row_pes_0_19_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_19_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_19_io_out_kv),
    .io_out_stage(global_row_pes_0_19_io_out_stage)
  );
  PE_1 global_row_pes_0_20 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_20_clock),
    .reset(global_row_pes_0_20_reset),
    .io_in_q(global_row_pes_0_20_io_in_q),
    .io_in_sum(global_row_pes_0_20_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_20_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_20_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_20_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_20_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_20_io_in_stage),
    .io_out_q(global_row_pes_0_20_io_out_q),
    .io_out_sum(global_row_pes_0_20_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_20_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_20_io_out_kv),
    .io_out_stage(global_row_pes_0_20_io_out_stage)
  );
  PE_1 global_row_pes_0_21 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_21_clock),
    .reset(global_row_pes_0_21_reset),
    .io_in_q(global_row_pes_0_21_io_in_q),
    .io_in_sum(global_row_pes_0_21_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_21_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_21_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_21_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_21_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_21_io_in_stage),
    .io_out_q(global_row_pes_0_21_io_out_q),
    .io_out_sum(global_row_pes_0_21_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_21_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_21_io_out_kv),
    .io_out_stage(global_row_pes_0_21_io_out_stage)
  );
  PE_1 global_row_pes_0_22 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_22_clock),
    .reset(global_row_pes_0_22_reset),
    .io_in_q(global_row_pes_0_22_io_in_q),
    .io_in_sum(global_row_pes_0_22_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_22_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_22_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_22_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_22_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_22_io_in_stage),
    .io_out_q(global_row_pes_0_22_io_out_q),
    .io_out_sum(global_row_pes_0_22_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_22_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_22_io_out_kv),
    .io_out_stage(global_row_pes_0_22_io_out_stage)
  );
  PE_1 global_row_pes_0_23 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_23_clock),
    .reset(global_row_pes_0_23_reset),
    .io_in_q(global_row_pes_0_23_io_in_q),
    .io_in_sum(global_row_pes_0_23_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_23_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_23_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_23_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_23_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_23_io_in_stage),
    .io_out_q(global_row_pes_0_23_io_out_q),
    .io_out_sum(global_row_pes_0_23_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_23_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_23_io_out_kv),
    .io_out_stage(global_row_pes_0_23_io_out_stage)
  );
  PE_1 global_row_pes_0_24 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_24_clock),
    .reset(global_row_pes_0_24_reset),
    .io_in_q(global_row_pes_0_24_io_in_q),
    .io_in_sum(global_row_pes_0_24_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_24_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_24_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_24_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_24_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_24_io_in_stage),
    .io_out_q(global_row_pes_0_24_io_out_q),
    .io_out_sum(global_row_pes_0_24_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_24_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_24_io_out_kv),
    .io_out_stage(global_row_pes_0_24_io_out_stage)
  );
  PE_1 global_row_pes_0_25 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_25_clock),
    .reset(global_row_pes_0_25_reset),
    .io_in_q(global_row_pes_0_25_io_in_q),
    .io_in_sum(global_row_pes_0_25_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_25_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_25_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_25_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_25_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_25_io_in_stage),
    .io_out_q(global_row_pes_0_25_io_out_q),
    .io_out_sum(global_row_pes_0_25_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_25_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_25_io_out_kv),
    .io_out_stage(global_row_pes_0_25_io_out_stage)
  );
  PE_1 global_row_pes_0_26 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_26_clock),
    .reset(global_row_pes_0_26_reset),
    .io_in_q(global_row_pes_0_26_io_in_q),
    .io_in_sum(global_row_pes_0_26_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_26_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_26_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_26_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_26_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_26_io_in_stage),
    .io_out_q(global_row_pes_0_26_io_out_q),
    .io_out_sum(global_row_pes_0_26_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_26_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_26_io_out_kv),
    .io_out_stage(global_row_pes_0_26_io_out_stage)
  );
  PE_1 global_row_pes_0_27 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_27_clock),
    .reset(global_row_pes_0_27_reset),
    .io_in_q(global_row_pes_0_27_io_in_q),
    .io_in_sum(global_row_pes_0_27_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_27_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_27_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_27_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_27_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_27_io_in_stage),
    .io_out_q(global_row_pes_0_27_io_out_q),
    .io_out_sum(global_row_pes_0_27_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_27_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_27_io_out_kv),
    .io_out_stage(global_row_pes_0_27_io_out_stage)
  );
  PE_1 global_row_pes_0_28 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_28_clock),
    .reset(global_row_pes_0_28_reset),
    .io_in_q(global_row_pes_0_28_io_in_q),
    .io_in_sum(global_row_pes_0_28_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_28_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_28_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_28_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_28_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_28_io_in_stage),
    .io_out_q(global_row_pes_0_28_io_out_q),
    .io_out_sum(global_row_pes_0_28_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_28_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_28_io_out_kv),
    .io_out_stage(global_row_pes_0_28_io_out_stage)
  );
  PE_1 global_row_pes_0_29 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_29_clock),
    .reset(global_row_pes_0_29_reset),
    .io_in_q(global_row_pes_0_29_io_in_q),
    .io_in_sum(global_row_pes_0_29_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_29_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_29_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_29_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_29_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_29_io_in_stage),
    .io_out_q(global_row_pes_0_29_io_out_q),
    .io_out_sum(global_row_pes_0_29_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_29_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_29_io_out_kv),
    .io_out_stage(global_row_pes_0_29_io_out_stage)
  );
  PE_1 global_row_pes_0_30 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_30_clock),
    .reset(global_row_pes_0_30_reset),
    .io_in_q(global_row_pes_0_30_io_in_q),
    .io_in_sum(global_row_pes_0_30_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_30_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_30_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_30_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_30_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_30_io_in_stage),
    .io_out_q(global_row_pes_0_30_io_out_q),
    .io_out_sum(global_row_pes_0_30_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_30_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_30_io_out_kv),
    .io_out_stage(global_row_pes_0_30_io_out_stage)
  );
  PE_1 global_row_pes_0_31 ( // @[PEArray.scala 29:49]
    .clock(global_row_pes_0_31_clock),
    .reset(global_row_pes_0_31_reset),
    .io_in_q(global_row_pes_0_31_io_in_q),
    .io_in_sum(global_row_pes_0_31_io_in_sum),
    .io_in_sum_exp(global_row_pes_0_31_io_in_sum_exp),
    .io_in_kv(global_row_pes_0_31_io_in_kv),
    .io_in_inv_sum_exp(global_row_pes_0_31_io_in_inv_sum_exp),
    .io_in_inv_sum(global_row_pes_0_31_io_in_inv_sum),
    .io_in_stage(global_row_pes_0_31_io_in_stage),
    .io_out_q(global_row_pes_0_31_io_out_q),
    .io_out_sum(global_row_pes_0_31_io_out_sum),
    .io_out_sum_exp(global_row_pes_0_31_io_out_sum_exp),
    .io_out_kv(global_row_pes_0_31_io_out_kv),
    .io_out_stage(global_row_pes_0_31_io_out_stage)
  );
  InverseModule inv_modules_0 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_0_io_in_sum),
    .io_in_exp(inv_modules_0_io_in_exp),
    .io_out_inv_sum(inv_modules_0_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_0_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_1 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_1_io_in_sum),
    .io_in_exp(inv_modules_1_io_in_exp),
    .io_out_inv_sum(inv_modules_1_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_1_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_2 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_2_io_in_sum),
    .io_in_exp(inv_modules_2_io_in_exp),
    .io_out_inv_sum(inv_modules_2_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_2_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_3 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_3_io_in_sum),
    .io_in_exp(inv_modules_3_io_in_exp),
    .io_out_inv_sum(inv_modules_3_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_3_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_4 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_4_io_in_sum),
    .io_in_exp(inv_modules_4_io_in_exp),
    .io_out_inv_sum(inv_modules_4_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_4_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_5 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_5_io_in_sum),
    .io_in_exp(inv_modules_5_io_in_exp),
    .io_out_inv_sum(inv_modules_5_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_5_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_6 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_6_io_in_sum),
    .io_in_exp(inv_modules_6_io_in_exp),
    .io_out_inv_sum(inv_modules_6_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_6_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_7 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_7_io_in_sum),
    .io_in_exp(inv_modules_7_io_in_exp),
    .io_out_inv_sum(inv_modules_7_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_7_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_8 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_8_io_in_sum),
    .io_in_exp(inv_modules_8_io_in_exp),
    .io_out_inv_sum(inv_modules_8_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_8_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_9 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_9_io_in_sum),
    .io_in_exp(inv_modules_9_io_in_exp),
    .io_out_inv_sum(inv_modules_9_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_9_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_10 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_10_io_in_sum),
    .io_in_exp(inv_modules_10_io_in_exp),
    .io_out_inv_sum(inv_modules_10_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_10_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_11 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_11_io_in_sum),
    .io_in_exp(inv_modules_11_io_in_exp),
    .io_out_inv_sum(inv_modules_11_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_11_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_12 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_12_io_in_sum),
    .io_in_exp(inv_modules_12_io_in_exp),
    .io_out_inv_sum(inv_modules_12_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_12_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_13 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_13_io_in_sum),
    .io_in_exp(inv_modules_13_io_in_exp),
    .io_out_inv_sum(inv_modules_13_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_13_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_14 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_14_io_in_sum),
    .io_in_exp(inv_modules_14_io_in_exp),
    .io_out_inv_sum(inv_modules_14_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_14_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_15 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_15_io_in_sum),
    .io_in_exp(inv_modules_15_io_in_exp),
    .io_out_inv_sum(inv_modules_15_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_15_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_16 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_16_io_in_sum),
    .io_in_exp(inv_modules_16_io_in_exp),
    .io_out_inv_sum(inv_modules_16_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_16_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_17 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_17_io_in_sum),
    .io_in_exp(inv_modules_17_io_in_exp),
    .io_out_inv_sum(inv_modules_17_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_17_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_18 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_18_io_in_sum),
    .io_in_exp(inv_modules_18_io_in_exp),
    .io_out_inv_sum(inv_modules_18_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_18_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_19 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_19_io_in_sum),
    .io_in_exp(inv_modules_19_io_in_exp),
    .io_out_inv_sum(inv_modules_19_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_19_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_20 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_20_io_in_sum),
    .io_in_exp(inv_modules_20_io_in_exp),
    .io_out_inv_sum(inv_modules_20_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_20_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_21 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_21_io_in_sum),
    .io_in_exp(inv_modules_21_io_in_exp),
    .io_out_inv_sum(inv_modules_21_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_21_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_22 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_22_io_in_sum),
    .io_in_exp(inv_modules_22_io_in_exp),
    .io_out_inv_sum(inv_modules_22_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_22_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_23 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_23_io_in_sum),
    .io_in_exp(inv_modules_23_io_in_exp),
    .io_out_inv_sum(inv_modules_23_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_23_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_24 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_24_io_in_sum),
    .io_in_exp(inv_modules_24_io_in_exp),
    .io_out_inv_sum(inv_modules_24_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_24_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_25 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_25_io_in_sum),
    .io_in_exp(inv_modules_25_io_in_exp),
    .io_out_inv_sum(inv_modules_25_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_25_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_26 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_26_io_in_sum),
    .io_in_exp(inv_modules_26_io_in_exp),
    .io_out_inv_sum(inv_modules_26_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_26_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_27 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_27_io_in_sum),
    .io_in_exp(inv_modules_27_io_in_exp),
    .io_out_inv_sum(inv_modules_27_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_27_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_28 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_28_io_in_sum),
    .io_in_exp(inv_modules_28_io_in_exp),
    .io_out_inv_sum(inv_modules_28_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_28_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_29 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_29_io_in_sum),
    .io_in_exp(inv_modules_29_io_in_exp),
    .io_out_inv_sum(inv_modules_29_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_29_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_30 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_30_io_in_sum),
    .io_in_exp(inv_modules_30_io_in_exp),
    .io_out_inv_sum(inv_modules_30_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_30_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_31 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_31_io_in_sum),
    .io_in_exp(inv_modules_31_io_in_exp),
    .io_out_inv_sum(inv_modules_31_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_31_io_out_inv_sum_exp)
  );
  InverseModule inv_modules_32 ( // @[PEArray.scala 31:73]
    .io_in_sum(inv_modules_32_io_in_sum),
    .io_in_exp(inv_modules_32_io_in_exp),
    .io_out_inv_sum(inv_modules_32_io_out_inv_sum),
    .io_out_inv_sum_exp(inv_modules_32_io_out_inv_sum_exp)
  );
  WeightedSumModule weighted_sum_modules_0 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_0_clock),
    .reset(weighted_sum_modules_0_reset),
    .io_in_sum(weighted_sum_modules_0_io_in_sum),
    .io_in_exp(weighted_sum_modules_0_io_in_exp),
    .io_control(weighted_sum_modules_0_io_control),
    .io_out_port(weighted_sum_modules_0_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_1 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_1_clock),
    .reset(weighted_sum_modules_1_reset),
    .io_in_sum(weighted_sum_modules_1_io_in_sum),
    .io_in_exp(weighted_sum_modules_1_io_in_exp),
    .io_control(weighted_sum_modules_1_io_control),
    .io_out_port(weighted_sum_modules_1_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_2 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_2_clock),
    .reset(weighted_sum_modules_2_reset),
    .io_in_sum(weighted_sum_modules_2_io_in_sum),
    .io_in_exp(weighted_sum_modules_2_io_in_exp),
    .io_control(weighted_sum_modules_2_io_control),
    .io_out_port(weighted_sum_modules_2_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_3 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_3_clock),
    .reset(weighted_sum_modules_3_reset),
    .io_in_sum(weighted_sum_modules_3_io_in_sum),
    .io_in_exp(weighted_sum_modules_3_io_in_exp),
    .io_control(weighted_sum_modules_3_io_control),
    .io_out_port(weighted_sum_modules_3_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_4 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_4_clock),
    .reset(weighted_sum_modules_4_reset),
    .io_in_sum(weighted_sum_modules_4_io_in_sum),
    .io_in_exp(weighted_sum_modules_4_io_in_exp),
    .io_control(weighted_sum_modules_4_io_control),
    .io_out_port(weighted_sum_modules_4_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_5 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_5_clock),
    .reset(weighted_sum_modules_5_reset),
    .io_in_sum(weighted_sum_modules_5_io_in_sum),
    .io_in_exp(weighted_sum_modules_5_io_in_exp),
    .io_control(weighted_sum_modules_5_io_control),
    .io_out_port(weighted_sum_modules_5_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_6 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_6_clock),
    .reset(weighted_sum_modules_6_reset),
    .io_in_sum(weighted_sum_modules_6_io_in_sum),
    .io_in_exp(weighted_sum_modules_6_io_in_exp),
    .io_control(weighted_sum_modules_6_io_control),
    .io_out_port(weighted_sum_modules_6_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_7 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_7_clock),
    .reset(weighted_sum_modules_7_reset),
    .io_in_sum(weighted_sum_modules_7_io_in_sum),
    .io_in_exp(weighted_sum_modules_7_io_in_exp),
    .io_control(weighted_sum_modules_7_io_control),
    .io_out_port(weighted_sum_modules_7_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_8 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_8_clock),
    .reset(weighted_sum_modules_8_reset),
    .io_in_sum(weighted_sum_modules_8_io_in_sum),
    .io_in_exp(weighted_sum_modules_8_io_in_exp),
    .io_control(weighted_sum_modules_8_io_control),
    .io_out_port(weighted_sum_modules_8_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_9 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_9_clock),
    .reset(weighted_sum_modules_9_reset),
    .io_in_sum(weighted_sum_modules_9_io_in_sum),
    .io_in_exp(weighted_sum_modules_9_io_in_exp),
    .io_control(weighted_sum_modules_9_io_control),
    .io_out_port(weighted_sum_modules_9_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_10 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_10_clock),
    .reset(weighted_sum_modules_10_reset),
    .io_in_sum(weighted_sum_modules_10_io_in_sum),
    .io_in_exp(weighted_sum_modules_10_io_in_exp),
    .io_control(weighted_sum_modules_10_io_control),
    .io_out_port(weighted_sum_modules_10_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_11 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_11_clock),
    .reset(weighted_sum_modules_11_reset),
    .io_in_sum(weighted_sum_modules_11_io_in_sum),
    .io_in_exp(weighted_sum_modules_11_io_in_exp),
    .io_control(weighted_sum_modules_11_io_control),
    .io_out_port(weighted_sum_modules_11_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_12 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_12_clock),
    .reset(weighted_sum_modules_12_reset),
    .io_in_sum(weighted_sum_modules_12_io_in_sum),
    .io_in_exp(weighted_sum_modules_12_io_in_exp),
    .io_control(weighted_sum_modules_12_io_control),
    .io_out_port(weighted_sum_modules_12_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_13 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_13_clock),
    .reset(weighted_sum_modules_13_reset),
    .io_in_sum(weighted_sum_modules_13_io_in_sum),
    .io_in_exp(weighted_sum_modules_13_io_in_exp),
    .io_control(weighted_sum_modules_13_io_control),
    .io_out_port(weighted_sum_modules_13_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_14 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_14_clock),
    .reset(weighted_sum_modules_14_reset),
    .io_in_sum(weighted_sum_modules_14_io_in_sum),
    .io_in_exp(weighted_sum_modules_14_io_in_exp),
    .io_control(weighted_sum_modules_14_io_control),
    .io_out_port(weighted_sum_modules_14_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_15 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_15_clock),
    .reset(weighted_sum_modules_15_reset),
    .io_in_sum(weighted_sum_modules_15_io_in_sum),
    .io_in_exp(weighted_sum_modules_15_io_in_exp),
    .io_control(weighted_sum_modules_15_io_control),
    .io_out_port(weighted_sum_modules_15_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_16 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_16_clock),
    .reset(weighted_sum_modules_16_reset),
    .io_in_sum(weighted_sum_modules_16_io_in_sum),
    .io_in_exp(weighted_sum_modules_16_io_in_exp),
    .io_control(weighted_sum_modules_16_io_control),
    .io_out_port(weighted_sum_modules_16_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_17 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_17_clock),
    .reset(weighted_sum_modules_17_reset),
    .io_in_sum(weighted_sum_modules_17_io_in_sum),
    .io_in_exp(weighted_sum_modules_17_io_in_exp),
    .io_control(weighted_sum_modules_17_io_control),
    .io_out_port(weighted_sum_modules_17_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_18 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_18_clock),
    .reset(weighted_sum_modules_18_reset),
    .io_in_sum(weighted_sum_modules_18_io_in_sum),
    .io_in_exp(weighted_sum_modules_18_io_in_exp),
    .io_control(weighted_sum_modules_18_io_control),
    .io_out_port(weighted_sum_modules_18_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_19 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_19_clock),
    .reset(weighted_sum_modules_19_reset),
    .io_in_sum(weighted_sum_modules_19_io_in_sum),
    .io_in_exp(weighted_sum_modules_19_io_in_exp),
    .io_control(weighted_sum_modules_19_io_control),
    .io_out_port(weighted_sum_modules_19_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_20 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_20_clock),
    .reset(weighted_sum_modules_20_reset),
    .io_in_sum(weighted_sum_modules_20_io_in_sum),
    .io_in_exp(weighted_sum_modules_20_io_in_exp),
    .io_control(weighted_sum_modules_20_io_control),
    .io_out_port(weighted_sum_modules_20_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_21 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_21_clock),
    .reset(weighted_sum_modules_21_reset),
    .io_in_sum(weighted_sum_modules_21_io_in_sum),
    .io_in_exp(weighted_sum_modules_21_io_in_exp),
    .io_control(weighted_sum_modules_21_io_control),
    .io_out_port(weighted_sum_modules_21_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_22 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_22_clock),
    .reset(weighted_sum_modules_22_reset),
    .io_in_sum(weighted_sum_modules_22_io_in_sum),
    .io_in_exp(weighted_sum_modules_22_io_in_exp),
    .io_control(weighted_sum_modules_22_io_control),
    .io_out_port(weighted_sum_modules_22_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_23 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_23_clock),
    .reset(weighted_sum_modules_23_reset),
    .io_in_sum(weighted_sum_modules_23_io_in_sum),
    .io_in_exp(weighted_sum_modules_23_io_in_exp),
    .io_control(weighted_sum_modules_23_io_control),
    .io_out_port(weighted_sum_modules_23_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_24 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_24_clock),
    .reset(weighted_sum_modules_24_reset),
    .io_in_sum(weighted_sum_modules_24_io_in_sum),
    .io_in_exp(weighted_sum_modules_24_io_in_exp),
    .io_control(weighted_sum_modules_24_io_control),
    .io_out_port(weighted_sum_modules_24_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_25 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_25_clock),
    .reset(weighted_sum_modules_25_reset),
    .io_in_sum(weighted_sum_modules_25_io_in_sum),
    .io_in_exp(weighted_sum_modules_25_io_in_exp),
    .io_control(weighted_sum_modules_25_io_control),
    .io_out_port(weighted_sum_modules_25_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_26 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_26_clock),
    .reset(weighted_sum_modules_26_reset),
    .io_in_sum(weighted_sum_modules_26_io_in_sum),
    .io_in_exp(weighted_sum_modules_26_io_in_exp),
    .io_control(weighted_sum_modules_26_io_control),
    .io_out_port(weighted_sum_modules_26_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_27 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_27_clock),
    .reset(weighted_sum_modules_27_reset),
    .io_in_sum(weighted_sum_modules_27_io_in_sum),
    .io_in_exp(weighted_sum_modules_27_io_in_exp),
    .io_control(weighted_sum_modules_27_io_control),
    .io_out_port(weighted_sum_modules_27_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_28 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_28_clock),
    .reset(weighted_sum_modules_28_reset),
    .io_in_sum(weighted_sum_modules_28_io_in_sum),
    .io_in_exp(weighted_sum_modules_28_io_in_exp),
    .io_control(weighted_sum_modules_28_io_control),
    .io_out_port(weighted_sum_modules_28_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_29 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_29_clock),
    .reset(weighted_sum_modules_29_reset),
    .io_in_sum(weighted_sum_modules_29_io_in_sum),
    .io_in_exp(weighted_sum_modules_29_io_in_exp),
    .io_control(weighted_sum_modules_29_io_control),
    .io_out_port(weighted_sum_modules_29_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_30 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_30_clock),
    .reset(weighted_sum_modules_30_reset),
    .io_in_sum(weighted_sum_modules_30_io_in_sum),
    .io_in_exp(weighted_sum_modules_30_io_in_exp),
    .io_control(weighted_sum_modules_30_io_control),
    .io_out_port(weighted_sum_modules_30_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_31 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_31_clock),
    .reset(weighted_sum_modules_31_reset),
    .io_in_sum(weighted_sum_modules_31_io_in_sum),
    .io_in_exp(weighted_sum_modules_31_io_in_exp),
    .io_control(weighted_sum_modules_31_io_control),
    .io_out_port(weighted_sum_modules_31_io_out_port)
  );
  WeightedSumModule weighted_sum_modules_32 ( // @[PEArray.scala 33:82]
    .clock(weighted_sum_modules_32_clock),
    .reset(weighted_sum_modules_32_reset),
    .io_in_sum(weighted_sum_modules_32_io_in_sum),
    .io_in_exp(weighted_sum_modules_32_io_in_exp),
    .io_control(weighted_sum_modules_32_io_control),
    .io_out_port(weighted_sum_modules_32_io_out_port)
  );
  assign io_out_ports_0 = weighted_sum_modules_0_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_1 = weighted_sum_modules_1_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_2 = weighted_sum_modules_2_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_3 = weighted_sum_modules_3_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_4 = weighted_sum_modules_4_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_5 = weighted_sum_modules_5_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_6 = weighted_sum_modules_6_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_7 = weighted_sum_modules_7_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_8 = weighted_sum_modules_8_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_9 = weighted_sum_modules_9_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_10 = weighted_sum_modules_10_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_11 = weighted_sum_modules_11_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_12 = weighted_sum_modules_12_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_13 = weighted_sum_modules_13_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_14 = weighted_sum_modules_14_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_15 = weighted_sum_modules_15_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_16 = weighted_sum_modules_16_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_17 = weighted_sum_modules_17_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_18 = weighted_sum_modules_18_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_19 = weighted_sum_modules_19_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_20 = weighted_sum_modules_20_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_21 = weighted_sum_modules_21_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_22 = weighted_sum_modules_22_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_23 = weighted_sum_modules_23_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_24 = weighted_sum_modules_24_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_25 = weighted_sum_modules_25_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_26 = weighted_sum_modules_26_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_27 = weighted_sum_modules_27_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_28 = weighted_sum_modules_28_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_29 = weighted_sum_modules_29_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_30 = weighted_sum_modules_30_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_31 = weighted_sum_modules_31_io_out_port; // @[PEArray.scala 98:25]
  assign io_out_ports_32 = weighted_sum_modules_32_io_out_port; // @[PEArray.scala 105:34]
  assign local_pes_0_0_clock = clock;
  assign local_pes_0_0_reset = reset;
  assign local_pes_0_0_io_in_q = io_q_ports_0; // @[PEArray.scala 51:37]
  assign local_pes_0_0_io_in_kv = io_kv_ports_31; // @[PEArray.scala 36:45]
  assign local_pes_0_0_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_0_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_0_io_in_stage = io_stage_ports_0; // @[PEArray.scala 52:41]
  assign local_pes_0_1_clock = clock;
  assign local_pes_0_1_reset = reset;
  assign local_pes_0_1_io_in_q = local_pes_0_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_1_io_in_sum = local_pes_0_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_0_1_io_in_kv = io_kv_ports_30; // @[PEArray.scala 36:45]
  assign local_pes_0_1_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_1_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_1_io_in_stage = local_pes_0_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_2_clock = clock;
  assign local_pes_0_2_reset = reset;
  assign local_pes_0_2_io_in_q = local_pes_0_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_2_io_in_sum = local_pes_0_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_2_io_in_sum_exp = local_pes_0_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_2_io_in_kv = io_kv_ports_29; // @[PEArray.scala 36:45]
  assign local_pes_0_2_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_2_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_2_io_in_stage = local_pes_0_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_3_clock = clock;
  assign local_pes_0_3_reset = reset;
  assign local_pes_0_3_io_in_q = local_pes_0_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_3_io_in_sum = local_pes_0_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_3_io_in_sum_exp = local_pes_0_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_3_io_in_kv = io_kv_ports_28; // @[PEArray.scala 36:45]
  assign local_pes_0_3_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_3_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_3_io_in_stage = local_pes_0_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_4_clock = clock;
  assign local_pes_0_4_reset = reset;
  assign local_pes_0_4_io_in_q = local_pes_0_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_4_io_in_sum = local_pes_0_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_4_io_in_sum_exp = local_pes_0_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_4_io_in_kv = io_kv_ports_27; // @[PEArray.scala 36:45]
  assign local_pes_0_4_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_4_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_4_io_in_stage = local_pes_0_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_5_clock = clock;
  assign local_pes_0_5_reset = reset;
  assign local_pes_0_5_io_in_q = local_pes_0_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_5_io_in_sum = local_pes_0_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_5_io_in_sum_exp = local_pes_0_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_5_io_in_kv = io_kv_ports_26; // @[PEArray.scala 36:45]
  assign local_pes_0_5_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_5_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_5_io_in_stage = local_pes_0_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_6_clock = clock;
  assign local_pes_0_6_reset = reset;
  assign local_pes_0_6_io_in_q = local_pes_0_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_6_io_in_sum = local_pes_0_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_6_io_in_sum_exp = local_pes_0_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_6_io_in_kv = io_kv_ports_25; // @[PEArray.scala 36:45]
  assign local_pes_0_6_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_6_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_6_io_in_stage = local_pes_0_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_7_clock = clock;
  assign local_pes_0_7_reset = reset;
  assign local_pes_0_7_io_in_q = local_pes_0_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_7_io_in_sum = local_pes_0_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_7_io_in_sum_exp = local_pes_0_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_7_io_in_kv = io_kv_ports_24; // @[PEArray.scala 36:45]
  assign local_pes_0_7_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_7_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_7_io_in_stage = local_pes_0_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_8_clock = clock;
  assign local_pes_0_8_reset = reset;
  assign local_pes_0_8_io_in_q = local_pes_0_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_8_io_in_sum = local_pes_0_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_8_io_in_sum_exp = local_pes_0_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_8_io_in_kv = io_kv_ports_23; // @[PEArray.scala 36:45]
  assign local_pes_0_8_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_8_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_8_io_in_stage = local_pes_0_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_9_clock = clock;
  assign local_pes_0_9_reset = reset;
  assign local_pes_0_9_io_in_q = local_pes_0_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_9_io_in_sum = local_pes_0_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_9_io_in_sum_exp = local_pes_0_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_9_io_in_kv = io_kv_ports_22; // @[PEArray.scala 36:45]
  assign local_pes_0_9_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_9_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_9_io_in_stage = local_pes_0_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_10_clock = clock;
  assign local_pes_0_10_reset = reset;
  assign local_pes_0_10_io_in_q = local_pes_0_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_10_io_in_sum = local_pes_0_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_10_io_in_sum_exp = local_pes_0_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_10_io_in_kv = io_kv_ports_21; // @[PEArray.scala 36:45]
  assign local_pes_0_10_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_10_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_10_io_in_stage = local_pes_0_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_11_clock = clock;
  assign local_pes_0_11_reset = reset;
  assign local_pes_0_11_io_in_q = local_pes_0_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_11_io_in_sum = local_pes_0_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_11_io_in_sum_exp = local_pes_0_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_11_io_in_kv = io_kv_ports_20; // @[PEArray.scala 36:45]
  assign local_pes_0_11_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_11_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_11_io_in_stage = local_pes_0_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_12_clock = clock;
  assign local_pes_0_12_reset = reset;
  assign local_pes_0_12_io_in_q = local_pes_0_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_12_io_in_sum = local_pes_0_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_12_io_in_sum_exp = local_pes_0_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_12_io_in_kv = io_kv_ports_19; // @[PEArray.scala 36:45]
  assign local_pes_0_12_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_12_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_12_io_in_stage = local_pes_0_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_13_clock = clock;
  assign local_pes_0_13_reset = reset;
  assign local_pes_0_13_io_in_q = local_pes_0_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_13_io_in_sum = local_pes_0_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_13_io_in_sum_exp = local_pes_0_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_13_io_in_kv = io_kv_ports_18; // @[PEArray.scala 36:45]
  assign local_pes_0_13_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_13_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_13_io_in_stage = local_pes_0_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_14_clock = clock;
  assign local_pes_0_14_reset = reset;
  assign local_pes_0_14_io_in_q = local_pes_0_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_14_io_in_sum = local_pes_0_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_14_io_in_sum_exp = local_pes_0_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_14_io_in_kv = io_kv_ports_17; // @[PEArray.scala 36:45]
  assign local_pes_0_14_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_14_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_14_io_in_stage = local_pes_0_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_15_clock = clock;
  assign local_pes_0_15_reset = reset;
  assign local_pes_0_15_io_in_q = local_pes_0_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_15_io_in_sum = local_pes_0_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_15_io_in_sum_exp = local_pes_0_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_15_io_in_kv = io_kv_ports_16; // @[PEArray.scala 36:45]
  assign local_pes_0_15_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_15_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_15_io_in_stage = local_pes_0_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_16_clock = clock;
  assign local_pes_0_16_reset = reset;
  assign local_pes_0_16_io_in_q = local_pes_0_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_16_io_in_sum = local_pes_0_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_16_io_in_sum_exp = local_pes_0_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_16_io_in_kv = io_kv_ports_15; // @[PEArray.scala 36:45]
  assign local_pes_0_16_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_16_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_16_io_in_stage = local_pes_0_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_17_clock = clock;
  assign local_pes_0_17_reset = reset;
  assign local_pes_0_17_io_in_q = local_pes_0_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_17_io_in_sum = local_pes_0_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_17_io_in_sum_exp = local_pes_0_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_17_io_in_kv = io_kv_ports_14; // @[PEArray.scala 36:45]
  assign local_pes_0_17_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_17_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_17_io_in_stage = local_pes_0_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_18_clock = clock;
  assign local_pes_0_18_reset = reset;
  assign local_pes_0_18_io_in_q = local_pes_0_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_18_io_in_sum = local_pes_0_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_18_io_in_sum_exp = local_pes_0_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_18_io_in_kv = io_kv_ports_13; // @[PEArray.scala 36:45]
  assign local_pes_0_18_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_18_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_18_io_in_stage = local_pes_0_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_19_clock = clock;
  assign local_pes_0_19_reset = reset;
  assign local_pes_0_19_io_in_q = local_pes_0_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_19_io_in_sum = local_pes_0_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_19_io_in_sum_exp = local_pes_0_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_19_io_in_kv = io_kv_ports_12; // @[PEArray.scala 36:45]
  assign local_pes_0_19_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_19_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_19_io_in_stage = local_pes_0_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_20_clock = clock;
  assign local_pes_0_20_reset = reset;
  assign local_pes_0_20_io_in_q = local_pes_0_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_20_io_in_sum = local_pes_0_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_20_io_in_sum_exp = local_pes_0_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_20_io_in_kv = io_kv_ports_11; // @[PEArray.scala 36:45]
  assign local_pes_0_20_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_20_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_20_io_in_stage = local_pes_0_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_21_clock = clock;
  assign local_pes_0_21_reset = reset;
  assign local_pes_0_21_io_in_q = local_pes_0_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_21_io_in_sum = local_pes_0_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_21_io_in_sum_exp = local_pes_0_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_21_io_in_kv = io_kv_ports_10; // @[PEArray.scala 36:45]
  assign local_pes_0_21_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_21_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_21_io_in_stage = local_pes_0_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_22_clock = clock;
  assign local_pes_0_22_reset = reset;
  assign local_pes_0_22_io_in_q = local_pes_0_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_22_io_in_sum = local_pes_0_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_22_io_in_sum_exp = local_pes_0_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_22_io_in_kv = io_kv_ports_9; // @[PEArray.scala 36:45]
  assign local_pes_0_22_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_22_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_22_io_in_stage = local_pes_0_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_23_clock = clock;
  assign local_pes_0_23_reset = reset;
  assign local_pes_0_23_io_in_q = local_pes_0_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_23_io_in_sum = local_pes_0_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_23_io_in_sum_exp = local_pes_0_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_23_io_in_kv = io_kv_ports_8; // @[PEArray.scala 36:45]
  assign local_pes_0_23_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_23_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_23_io_in_stage = local_pes_0_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_24_clock = clock;
  assign local_pes_0_24_reset = reset;
  assign local_pes_0_24_io_in_q = local_pes_0_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_24_io_in_sum = local_pes_0_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_24_io_in_sum_exp = local_pes_0_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_24_io_in_kv = io_kv_ports_7; // @[PEArray.scala 36:45]
  assign local_pes_0_24_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_24_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_24_io_in_stage = local_pes_0_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_25_clock = clock;
  assign local_pes_0_25_reset = reset;
  assign local_pes_0_25_io_in_q = local_pes_0_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_25_io_in_sum = local_pes_0_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_25_io_in_sum_exp = local_pes_0_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_25_io_in_kv = io_kv_ports_6; // @[PEArray.scala 36:45]
  assign local_pes_0_25_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_25_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_25_io_in_stage = local_pes_0_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_26_clock = clock;
  assign local_pes_0_26_reset = reset;
  assign local_pes_0_26_io_in_q = local_pes_0_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_26_io_in_sum = local_pes_0_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_26_io_in_sum_exp = local_pes_0_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_26_io_in_kv = io_kv_ports_5; // @[PEArray.scala 36:45]
  assign local_pes_0_26_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_26_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_26_io_in_stage = local_pes_0_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_27_clock = clock;
  assign local_pes_0_27_reset = reset;
  assign local_pes_0_27_io_in_q = local_pes_0_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_27_io_in_sum = local_pes_0_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_27_io_in_sum_exp = local_pes_0_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_27_io_in_kv = io_kv_ports_4; // @[PEArray.scala 36:45]
  assign local_pes_0_27_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_27_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_27_io_in_stage = local_pes_0_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_28_clock = clock;
  assign local_pes_0_28_reset = reset;
  assign local_pes_0_28_io_in_q = local_pes_0_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_28_io_in_sum = local_pes_0_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_28_io_in_sum_exp = local_pes_0_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_28_io_in_kv = io_kv_ports_3; // @[PEArray.scala 36:45]
  assign local_pes_0_28_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_28_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_28_io_in_stage = local_pes_0_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_29_clock = clock;
  assign local_pes_0_29_reset = reset;
  assign local_pes_0_29_io_in_q = local_pes_0_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_29_io_in_sum = local_pes_0_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_29_io_in_sum_exp = local_pes_0_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_29_io_in_kv = io_kv_ports_2; // @[PEArray.scala 36:45]
  assign local_pes_0_29_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_29_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_29_io_in_stage = local_pes_0_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_30_clock = clock;
  assign local_pes_0_30_reset = reset;
  assign local_pes_0_30_io_in_q = local_pes_0_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_30_io_in_sum = local_pes_0_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_30_io_in_sum_exp = local_pes_0_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_30_io_in_kv = io_kv_ports_1; // @[PEArray.scala 36:45]
  assign local_pes_0_30_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_30_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_30_io_in_stage = local_pes_0_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_0_31_clock = clock;
  assign local_pes_0_31_reset = reset;
  assign local_pes_0_31_io_in_q = local_pes_0_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_0_31_io_in_sum = local_pes_0_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_0_31_io_in_sum_exp = local_pes_0_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_0_31_io_in_kv = io_kv_ports_0; // @[PEArray.scala 36:45]
  assign local_pes_0_31_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_0_31_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_0_31_io_in_stage = local_pes_0_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_0_clock = clock;
  assign local_pes_1_0_reset = reset;
  assign local_pes_1_0_io_in_q = io_q_ports_1; // @[PEArray.scala 51:37]
  assign local_pes_1_0_io_in_kv = io_kv_ports_32; // @[PEArray.scala 40:34]
  assign local_pes_1_0_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_0_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_0_io_in_stage = io_stage_ports_1; // @[PEArray.scala 52:41]
  assign local_pes_1_1_clock = clock;
  assign local_pes_1_1_reset = reset;
  assign local_pes_1_1_io_in_q = local_pes_1_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_1_io_in_sum = local_pes_1_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_1_1_io_in_kv = local_pes_0_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_1_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_1_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_1_io_in_stage = local_pes_1_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_2_clock = clock;
  assign local_pes_1_2_reset = reset;
  assign local_pes_1_2_io_in_q = local_pes_1_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_2_io_in_sum = local_pes_1_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_2_io_in_sum_exp = local_pes_1_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_2_io_in_kv = local_pes_0_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_2_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_2_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_2_io_in_stage = local_pes_1_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_3_clock = clock;
  assign local_pes_1_3_reset = reset;
  assign local_pes_1_3_io_in_q = local_pes_1_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_3_io_in_sum = local_pes_1_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_3_io_in_sum_exp = local_pes_1_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_3_io_in_kv = local_pes_0_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_3_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_3_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_3_io_in_stage = local_pes_1_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_4_clock = clock;
  assign local_pes_1_4_reset = reset;
  assign local_pes_1_4_io_in_q = local_pes_1_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_4_io_in_sum = local_pes_1_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_4_io_in_sum_exp = local_pes_1_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_4_io_in_kv = local_pes_0_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_4_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_4_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_4_io_in_stage = local_pes_1_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_5_clock = clock;
  assign local_pes_1_5_reset = reset;
  assign local_pes_1_5_io_in_q = local_pes_1_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_5_io_in_sum = local_pes_1_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_5_io_in_sum_exp = local_pes_1_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_5_io_in_kv = local_pes_0_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_5_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_5_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_5_io_in_stage = local_pes_1_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_6_clock = clock;
  assign local_pes_1_6_reset = reset;
  assign local_pes_1_6_io_in_q = local_pes_1_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_6_io_in_sum = local_pes_1_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_6_io_in_sum_exp = local_pes_1_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_6_io_in_kv = local_pes_0_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_6_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_6_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_6_io_in_stage = local_pes_1_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_7_clock = clock;
  assign local_pes_1_7_reset = reset;
  assign local_pes_1_7_io_in_q = local_pes_1_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_7_io_in_sum = local_pes_1_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_7_io_in_sum_exp = local_pes_1_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_7_io_in_kv = local_pes_0_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_7_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_7_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_7_io_in_stage = local_pes_1_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_8_clock = clock;
  assign local_pes_1_8_reset = reset;
  assign local_pes_1_8_io_in_q = local_pes_1_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_8_io_in_sum = local_pes_1_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_8_io_in_sum_exp = local_pes_1_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_8_io_in_kv = local_pes_0_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_8_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_8_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_8_io_in_stage = local_pes_1_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_9_clock = clock;
  assign local_pes_1_9_reset = reset;
  assign local_pes_1_9_io_in_q = local_pes_1_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_9_io_in_sum = local_pes_1_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_9_io_in_sum_exp = local_pes_1_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_9_io_in_kv = local_pes_0_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_9_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_9_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_9_io_in_stage = local_pes_1_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_10_clock = clock;
  assign local_pes_1_10_reset = reset;
  assign local_pes_1_10_io_in_q = local_pes_1_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_10_io_in_sum = local_pes_1_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_10_io_in_sum_exp = local_pes_1_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_10_io_in_kv = local_pes_0_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_10_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_10_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_10_io_in_stage = local_pes_1_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_11_clock = clock;
  assign local_pes_1_11_reset = reset;
  assign local_pes_1_11_io_in_q = local_pes_1_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_11_io_in_sum = local_pes_1_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_11_io_in_sum_exp = local_pes_1_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_11_io_in_kv = local_pes_0_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_11_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_11_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_11_io_in_stage = local_pes_1_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_12_clock = clock;
  assign local_pes_1_12_reset = reset;
  assign local_pes_1_12_io_in_q = local_pes_1_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_12_io_in_sum = local_pes_1_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_12_io_in_sum_exp = local_pes_1_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_12_io_in_kv = local_pes_0_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_12_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_12_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_12_io_in_stage = local_pes_1_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_13_clock = clock;
  assign local_pes_1_13_reset = reset;
  assign local_pes_1_13_io_in_q = local_pes_1_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_13_io_in_sum = local_pes_1_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_13_io_in_sum_exp = local_pes_1_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_13_io_in_kv = local_pes_0_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_13_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_13_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_13_io_in_stage = local_pes_1_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_14_clock = clock;
  assign local_pes_1_14_reset = reset;
  assign local_pes_1_14_io_in_q = local_pes_1_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_14_io_in_sum = local_pes_1_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_14_io_in_sum_exp = local_pes_1_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_14_io_in_kv = local_pes_0_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_14_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_14_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_14_io_in_stage = local_pes_1_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_15_clock = clock;
  assign local_pes_1_15_reset = reset;
  assign local_pes_1_15_io_in_q = local_pes_1_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_15_io_in_sum = local_pes_1_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_15_io_in_sum_exp = local_pes_1_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_15_io_in_kv = local_pes_0_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_15_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_15_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_15_io_in_stage = local_pes_1_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_16_clock = clock;
  assign local_pes_1_16_reset = reset;
  assign local_pes_1_16_io_in_q = local_pes_1_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_16_io_in_sum = local_pes_1_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_16_io_in_sum_exp = local_pes_1_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_16_io_in_kv = local_pes_0_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_16_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_16_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_16_io_in_stage = local_pes_1_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_17_clock = clock;
  assign local_pes_1_17_reset = reset;
  assign local_pes_1_17_io_in_q = local_pes_1_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_17_io_in_sum = local_pes_1_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_17_io_in_sum_exp = local_pes_1_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_17_io_in_kv = local_pes_0_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_17_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_17_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_17_io_in_stage = local_pes_1_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_18_clock = clock;
  assign local_pes_1_18_reset = reset;
  assign local_pes_1_18_io_in_q = local_pes_1_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_18_io_in_sum = local_pes_1_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_18_io_in_sum_exp = local_pes_1_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_18_io_in_kv = local_pes_0_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_18_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_18_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_18_io_in_stage = local_pes_1_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_19_clock = clock;
  assign local_pes_1_19_reset = reset;
  assign local_pes_1_19_io_in_q = local_pes_1_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_19_io_in_sum = local_pes_1_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_19_io_in_sum_exp = local_pes_1_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_19_io_in_kv = local_pes_0_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_19_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_19_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_19_io_in_stage = local_pes_1_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_20_clock = clock;
  assign local_pes_1_20_reset = reset;
  assign local_pes_1_20_io_in_q = local_pes_1_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_20_io_in_sum = local_pes_1_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_20_io_in_sum_exp = local_pes_1_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_20_io_in_kv = local_pes_0_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_20_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_20_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_20_io_in_stage = local_pes_1_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_21_clock = clock;
  assign local_pes_1_21_reset = reset;
  assign local_pes_1_21_io_in_q = local_pes_1_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_21_io_in_sum = local_pes_1_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_21_io_in_sum_exp = local_pes_1_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_21_io_in_kv = local_pes_0_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_21_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_21_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_21_io_in_stage = local_pes_1_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_22_clock = clock;
  assign local_pes_1_22_reset = reset;
  assign local_pes_1_22_io_in_q = local_pes_1_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_22_io_in_sum = local_pes_1_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_22_io_in_sum_exp = local_pes_1_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_22_io_in_kv = local_pes_0_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_22_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_22_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_22_io_in_stage = local_pes_1_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_23_clock = clock;
  assign local_pes_1_23_reset = reset;
  assign local_pes_1_23_io_in_q = local_pes_1_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_23_io_in_sum = local_pes_1_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_23_io_in_sum_exp = local_pes_1_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_23_io_in_kv = local_pes_0_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_23_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_23_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_23_io_in_stage = local_pes_1_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_24_clock = clock;
  assign local_pes_1_24_reset = reset;
  assign local_pes_1_24_io_in_q = local_pes_1_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_24_io_in_sum = local_pes_1_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_24_io_in_sum_exp = local_pes_1_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_24_io_in_kv = local_pes_0_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_24_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_24_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_24_io_in_stage = local_pes_1_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_25_clock = clock;
  assign local_pes_1_25_reset = reset;
  assign local_pes_1_25_io_in_q = local_pes_1_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_25_io_in_sum = local_pes_1_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_25_io_in_sum_exp = local_pes_1_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_25_io_in_kv = local_pes_0_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_25_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_25_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_25_io_in_stage = local_pes_1_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_26_clock = clock;
  assign local_pes_1_26_reset = reset;
  assign local_pes_1_26_io_in_q = local_pes_1_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_26_io_in_sum = local_pes_1_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_26_io_in_sum_exp = local_pes_1_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_26_io_in_kv = local_pes_0_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_26_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_26_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_26_io_in_stage = local_pes_1_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_27_clock = clock;
  assign local_pes_1_27_reset = reset;
  assign local_pes_1_27_io_in_q = local_pes_1_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_27_io_in_sum = local_pes_1_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_27_io_in_sum_exp = local_pes_1_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_27_io_in_kv = local_pes_0_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_27_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_27_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_27_io_in_stage = local_pes_1_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_28_clock = clock;
  assign local_pes_1_28_reset = reset;
  assign local_pes_1_28_io_in_q = local_pes_1_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_28_io_in_sum = local_pes_1_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_28_io_in_sum_exp = local_pes_1_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_28_io_in_kv = local_pes_0_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_28_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_28_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_28_io_in_stage = local_pes_1_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_29_clock = clock;
  assign local_pes_1_29_reset = reset;
  assign local_pes_1_29_io_in_q = local_pes_1_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_29_io_in_sum = local_pes_1_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_29_io_in_sum_exp = local_pes_1_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_29_io_in_kv = local_pes_0_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_29_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_29_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_29_io_in_stage = local_pes_1_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_30_clock = clock;
  assign local_pes_1_30_reset = reset;
  assign local_pes_1_30_io_in_q = local_pes_1_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_30_io_in_sum = local_pes_1_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_30_io_in_sum_exp = local_pes_1_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_30_io_in_kv = local_pes_0_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_30_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_30_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_30_io_in_stage = local_pes_1_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_1_31_clock = clock;
  assign local_pes_1_31_reset = reset;
  assign local_pes_1_31_io_in_q = local_pes_1_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_1_31_io_in_sum = local_pes_1_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_1_31_io_in_sum_exp = local_pes_1_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_1_31_io_in_kv = local_pes_0_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_1_31_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_1_31_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_1_31_io_in_stage = local_pes_1_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_0_clock = clock;
  assign local_pes_2_0_reset = reset;
  assign local_pes_2_0_io_in_q = io_q_ports_2; // @[PEArray.scala 51:37]
  assign local_pes_2_0_io_in_kv = io_kv_ports_33; // @[PEArray.scala 40:34]
  assign local_pes_2_0_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_0_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_0_io_in_stage = io_stage_ports_2; // @[PEArray.scala 52:41]
  assign local_pes_2_1_clock = clock;
  assign local_pes_2_1_reset = reset;
  assign local_pes_2_1_io_in_q = local_pes_2_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_1_io_in_sum = local_pes_2_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_2_1_io_in_kv = local_pes_1_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_1_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_1_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_1_io_in_stage = local_pes_2_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_2_clock = clock;
  assign local_pes_2_2_reset = reset;
  assign local_pes_2_2_io_in_q = local_pes_2_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_2_io_in_sum = local_pes_2_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_2_io_in_sum_exp = local_pes_2_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_2_io_in_kv = local_pes_1_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_2_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_2_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_2_io_in_stage = local_pes_2_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_3_clock = clock;
  assign local_pes_2_3_reset = reset;
  assign local_pes_2_3_io_in_q = local_pes_2_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_3_io_in_sum = local_pes_2_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_3_io_in_sum_exp = local_pes_2_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_3_io_in_kv = local_pes_1_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_3_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_3_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_3_io_in_stage = local_pes_2_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_4_clock = clock;
  assign local_pes_2_4_reset = reset;
  assign local_pes_2_4_io_in_q = local_pes_2_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_4_io_in_sum = local_pes_2_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_4_io_in_sum_exp = local_pes_2_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_4_io_in_kv = local_pes_1_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_4_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_4_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_4_io_in_stage = local_pes_2_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_5_clock = clock;
  assign local_pes_2_5_reset = reset;
  assign local_pes_2_5_io_in_q = local_pes_2_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_5_io_in_sum = local_pes_2_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_5_io_in_sum_exp = local_pes_2_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_5_io_in_kv = local_pes_1_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_5_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_5_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_5_io_in_stage = local_pes_2_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_6_clock = clock;
  assign local_pes_2_6_reset = reset;
  assign local_pes_2_6_io_in_q = local_pes_2_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_6_io_in_sum = local_pes_2_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_6_io_in_sum_exp = local_pes_2_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_6_io_in_kv = local_pes_1_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_6_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_6_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_6_io_in_stage = local_pes_2_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_7_clock = clock;
  assign local_pes_2_7_reset = reset;
  assign local_pes_2_7_io_in_q = local_pes_2_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_7_io_in_sum = local_pes_2_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_7_io_in_sum_exp = local_pes_2_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_7_io_in_kv = local_pes_1_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_7_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_7_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_7_io_in_stage = local_pes_2_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_8_clock = clock;
  assign local_pes_2_8_reset = reset;
  assign local_pes_2_8_io_in_q = local_pes_2_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_8_io_in_sum = local_pes_2_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_8_io_in_sum_exp = local_pes_2_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_8_io_in_kv = local_pes_1_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_8_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_8_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_8_io_in_stage = local_pes_2_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_9_clock = clock;
  assign local_pes_2_9_reset = reset;
  assign local_pes_2_9_io_in_q = local_pes_2_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_9_io_in_sum = local_pes_2_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_9_io_in_sum_exp = local_pes_2_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_9_io_in_kv = local_pes_1_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_9_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_9_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_9_io_in_stage = local_pes_2_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_10_clock = clock;
  assign local_pes_2_10_reset = reset;
  assign local_pes_2_10_io_in_q = local_pes_2_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_10_io_in_sum = local_pes_2_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_10_io_in_sum_exp = local_pes_2_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_10_io_in_kv = local_pes_1_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_10_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_10_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_10_io_in_stage = local_pes_2_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_11_clock = clock;
  assign local_pes_2_11_reset = reset;
  assign local_pes_2_11_io_in_q = local_pes_2_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_11_io_in_sum = local_pes_2_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_11_io_in_sum_exp = local_pes_2_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_11_io_in_kv = local_pes_1_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_11_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_11_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_11_io_in_stage = local_pes_2_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_12_clock = clock;
  assign local_pes_2_12_reset = reset;
  assign local_pes_2_12_io_in_q = local_pes_2_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_12_io_in_sum = local_pes_2_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_12_io_in_sum_exp = local_pes_2_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_12_io_in_kv = local_pes_1_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_12_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_12_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_12_io_in_stage = local_pes_2_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_13_clock = clock;
  assign local_pes_2_13_reset = reset;
  assign local_pes_2_13_io_in_q = local_pes_2_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_13_io_in_sum = local_pes_2_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_13_io_in_sum_exp = local_pes_2_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_13_io_in_kv = local_pes_1_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_13_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_13_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_13_io_in_stage = local_pes_2_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_14_clock = clock;
  assign local_pes_2_14_reset = reset;
  assign local_pes_2_14_io_in_q = local_pes_2_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_14_io_in_sum = local_pes_2_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_14_io_in_sum_exp = local_pes_2_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_14_io_in_kv = local_pes_1_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_14_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_14_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_14_io_in_stage = local_pes_2_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_15_clock = clock;
  assign local_pes_2_15_reset = reset;
  assign local_pes_2_15_io_in_q = local_pes_2_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_15_io_in_sum = local_pes_2_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_15_io_in_sum_exp = local_pes_2_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_15_io_in_kv = local_pes_1_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_15_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_15_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_15_io_in_stage = local_pes_2_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_16_clock = clock;
  assign local_pes_2_16_reset = reset;
  assign local_pes_2_16_io_in_q = local_pes_2_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_16_io_in_sum = local_pes_2_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_16_io_in_sum_exp = local_pes_2_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_16_io_in_kv = local_pes_1_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_16_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_16_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_16_io_in_stage = local_pes_2_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_17_clock = clock;
  assign local_pes_2_17_reset = reset;
  assign local_pes_2_17_io_in_q = local_pes_2_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_17_io_in_sum = local_pes_2_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_17_io_in_sum_exp = local_pes_2_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_17_io_in_kv = local_pes_1_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_17_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_17_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_17_io_in_stage = local_pes_2_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_18_clock = clock;
  assign local_pes_2_18_reset = reset;
  assign local_pes_2_18_io_in_q = local_pes_2_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_18_io_in_sum = local_pes_2_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_18_io_in_sum_exp = local_pes_2_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_18_io_in_kv = local_pes_1_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_18_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_18_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_18_io_in_stage = local_pes_2_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_19_clock = clock;
  assign local_pes_2_19_reset = reset;
  assign local_pes_2_19_io_in_q = local_pes_2_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_19_io_in_sum = local_pes_2_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_19_io_in_sum_exp = local_pes_2_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_19_io_in_kv = local_pes_1_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_19_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_19_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_19_io_in_stage = local_pes_2_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_20_clock = clock;
  assign local_pes_2_20_reset = reset;
  assign local_pes_2_20_io_in_q = local_pes_2_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_20_io_in_sum = local_pes_2_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_20_io_in_sum_exp = local_pes_2_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_20_io_in_kv = local_pes_1_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_20_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_20_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_20_io_in_stage = local_pes_2_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_21_clock = clock;
  assign local_pes_2_21_reset = reset;
  assign local_pes_2_21_io_in_q = local_pes_2_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_21_io_in_sum = local_pes_2_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_21_io_in_sum_exp = local_pes_2_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_21_io_in_kv = local_pes_1_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_21_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_21_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_21_io_in_stage = local_pes_2_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_22_clock = clock;
  assign local_pes_2_22_reset = reset;
  assign local_pes_2_22_io_in_q = local_pes_2_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_22_io_in_sum = local_pes_2_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_22_io_in_sum_exp = local_pes_2_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_22_io_in_kv = local_pes_1_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_22_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_22_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_22_io_in_stage = local_pes_2_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_23_clock = clock;
  assign local_pes_2_23_reset = reset;
  assign local_pes_2_23_io_in_q = local_pes_2_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_23_io_in_sum = local_pes_2_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_23_io_in_sum_exp = local_pes_2_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_23_io_in_kv = local_pes_1_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_23_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_23_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_23_io_in_stage = local_pes_2_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_24_clock = clock;
  assign local_pes_2_24_reset = reset;
  assign local_pes_2_24_io_in_q = local_pes_2_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_24_io_in_sum = local_pes_2_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_24_io_in_sum_exp = local_pes_2_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_24_io_in_kv = local_pes_1_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_24_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_24_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_24_io_in_stage = local_pes_2_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_25_clock = clock;
  assign local_pes_2_25_reset = reset;
  assign local_pes_2_25_io_in_q = local_pes_2_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_25_io_in_sum = local_pes_2_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_25_io_in_sum_exp = local_pes_2_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_25_io_in_kv = local_pes_1_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_25_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_25_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_25_io_in_stage = local_pes_2_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_26_clock = clock;
  assign local_pes_2_26_reset = reset;
  assign local_pes_2_26_io_in_q = local_pes_2_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_26_io_in_sum = local_pes_2_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_26_io_in_sum_exp = local_pes_2_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_26_io_in_kv = local_pes_1_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_26_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_26_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_26_io_in_stage = local_pes_2_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_27_clock = clock;
  assign local_pes_2_27_reset = reset;
  assign local_pes_2_27_io_in_q = local_pes_2_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_27_io_in_sum = local_pes_2_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_27_io_in_sum_exp = local_pes_2_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_27_io_in_kv = local_pes_1_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_27_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_27_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_27_io_in_stage = local_pes_2_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_28_clock = clock;
  assign local_pes_2_28_reset = reset;
  assign local_pes_2_28_io_in_q = local_pes_2_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_28_io_in_sum = local_pes_2_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_28_io_in_sum_exp = local_pes_2_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_28_io_in_kv = local_pes_1_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_28_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_28_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_28_io_in_stage = local_pes_2_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_29_clock = clock;
  assign local_pes_2_29_reset = reset;
  assign local_pes_2_29_io_in_q = local_pes_2_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_29_io_in_sum = local_pes_2_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_29_io_in_sum_exp = local_pes_2_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_29_io_in_kv = local_pes_1_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_29_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_29_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_29_io_in_stage = local_pes_2_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_30_clock = clock;
  assign local_pes_2_30_reset = reset;
  assign local_pes_2_30_io_in_q = local_pes_2_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_30_io_in_sum = local_pes_2_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_30_io_in_sum_exp = local_pes_2_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_30_io_in_kv = local_pes_1_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_30_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_30_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_30_io_in_stage = local_pes_2_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_2_31_clock = clock;
  assign local_pes_2_31_reset = reset;
  assign local_pes_2_31_io_in_q = local_pes_2_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_2_31_io_in_sum = local_pes_2_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_2_31_io_in_sum_exp = local_pes_2_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_2_31_io_in_kv = local_pes_1_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_2_31_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_2_31_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_2_31_io_in_stage = local_pes_2_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_0_clock = clock;
  assign local_pes_3_0_reset = reset;
  assign local_pes_3_0_io_in_q = io_q_ports_3; // @[PEArray.scala 51:37]
  assign local_pes_3_0_io_in_kv = io_kv_ports_34; // @[PEArray.scala 40:34]
  assign local_pes_3_0_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_0_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_0_io_in_stage = io_stage_ports_3; // @[PEArray.scala 52:41]
  assign local_pes_3_1_clock = clock;
  assign local_pes_3_1_reset = reset;
  assign local_pes_3_1_io_in_q = local_pes_3_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_1_io_in_sum = local_pes_3_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_3_1_io_in_kv = local_pes_2_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_1_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_1_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_1_io_in_stage = local_pes_3_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_2_clock = clock;
  assign local_pes_3_2_reset = reset;
  assign local_pes_3_2_io_in_q = local_pes_3_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_2_io_in_sum = local_pes_3_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_2_io_in_sum_exp = local_pes_3_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_2_io_in_kv = local_pes_2_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_2_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_2_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_2_io_in_stage = local_pes_3_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_3_clock = clock;
  assign local_pes_3_3_reset = reset;
  assign local_pes_3_3_io_in_q = local_pes_3_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_3_io_in_sum = local_pes_3_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_3_io_in_sum_exp = local_pes_3_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_3_io_in_kv = local_pes_2_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_3_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_3_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_3_io_in_stage = local_pes_3_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_4_clock = clock;
  assign local_pes_3_4_reset = reset;
  assign local_pes_3_4_io_in_q = local_pes_3_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_4_io_in_sum = local_pes_3_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_4_io_in_sum_exp = local_pes_3_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_4_io_in_kv = local_pes_2_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_4_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_4_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_4_io_in_stage = local_pes_3_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_5_clock = clock;
  assign local_pes_3_5_reset = reset;
  assign local_pes_3_5_io_in_q = local_pes_3_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_5_io_in_sum = local_pes_3_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_5_io_in_sum_exp = local_pes_3_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_5_io_in_kv = local_pes_2_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_5_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_5_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_5_io_in_stage = local_pes_3_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_6_clock = clock;
  assign local_pes_3_6_reset = reset;
  assign local_pes_3_6_io_in_q = local_pes_3_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_6_io_in_sum = local_pes_3_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_6_io_in_sum_exp = local_pes_3_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_6_io_in_kv = local_pes_2_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_6_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_6_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_6_io_in_stage = local_pes_3_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_7_clock = clock;
  assign local_pes_3_7_reset = reset;
  assign local_pes_3_7_io_in_q = local_pes_3_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_7_io_in_sum = local_pes_3_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_7_io_in_sum_exp = local_pes_3_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_7_io_in_kv = local_pes_2_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_7_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_7_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_7_io_in_stage = local_pes_3_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_8_clock = clock;
  assign local_pes_3_8_reset = reset;
  assign local_pes_3_8_io_in_q = local_pes_3_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_8_io_in_sum = local_pes_3_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_8_io_in_sum_exp = local_pes_3_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_8_io_in_kv = local_pes_2_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_8_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_8_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_8_io_in_stage = local_pes_3_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_9_clock = clock;
  assign local_pes_3_9_reset = reset;
  assign local_pes_3_9_io_in_q = local_pes_3_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_9_io_in_sum = local_pes_3_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_9_io_in_sum_exp = local_pes_3_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_9_io_in_kv = local_pes_2_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_9_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_9_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_9_io_in_stage = local_pes_3_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_10_clock = clock;
  assign local_pes_3_10_reset = reset;
  assign local_pes_3_10_io_in_q = local_pes_3_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_10_io_in_sum = local_pes_3_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_10_io_in_sum_exp = local_pes_3_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_10_io_in_kv = local_pes_2_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_10_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_10_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_10_io_in_stage = local_pes_3_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_11_clock = clock;
  assign local_pes_3_11_reset = reset;
  assign local_pes_3_11_io_in_q = local_pes_3_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_11_io_in_sum = local_pes_3_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_11_io_in_sum_exp = local_pes_3_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_11_io_in_kv = local_pes_2_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_11_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_11_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_11_io_in_stage = local_pes_3_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_12_clock = clock;
  assign local_pes_3_12_reset = reset;
  assign local_pes_3_12_io_in_q = local_pes_3_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_12_io_in_sum = local_pes_3_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_12_io_in_sum_exp = local_pes_3_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_12_io_in_kv = local_pes_2_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_12_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_12_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_12_io_in_stage = local_pes_3_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_13_clock = clock;
  assign local_pes_3_13_reset = reset;
  assign local_pes_3_13_io_in_q = local_pes_3_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_13_io_in_sum = local_pes_3_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_13_io_in_sum_exp = local_pes_3_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_13_io_in_kv = local_pes_2_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_13_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_13_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_13_io_in_stage = local_pes_3_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_14_clock = clock;
  assign local_pes_3_14_reset = reset;
  assign local_pes_3_14_io_in_q = local_pes_3_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_14_io_in_sum = local_pes_3_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_14_io_in_sum_exp = local_pes_3_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_14_io_in_kv = local_pes_2_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_14_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_14_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_14_io_in_stage = local_pes_3_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_15_clock = clock;
  assign local_pes_3_15_reset = reset;
  assign local_pes_3_15_io_in_q = local_pes_3_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_15_io_in_sum = local_pes_3_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_15_io_in_sum_exp = local_pes_3_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_15_io_in_kv = local_pes_2_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_15_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_15_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_15_io_in_stage = local_pes_3_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_16_clock = clock;
  assign local_pes_3_16_reset = reset;
  assign local_pes_3_16_io_in_q = local_pes_3_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_16_io_in_sum = local_pes_3_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_16_io_in_sum_exp = local_pes_3_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_16_io_in_kv = local_pes_2_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_16_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_16_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_16_io_in_stage = local_pes_3_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_17_clock = clock;
  assign local_pes_3_17_reset = reset;
  assign local_pes_3_17_io_in_q = local_pes_3_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_17_io_in_sum = local_pes_3_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_17_io_in_sum_exp = local_pes_3_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_17_io_in_kv = local_pes_2_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_17_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_17_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_17_io_in_stage = local_pes_3_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_18_clock = clock;
  assign local_pes_3_18_reset = reset;
  assign local_pes_3_18_io_in_q = local_pes_3_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_18_io_in_sum = local_pes_3_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_18_io_in_sum_exp = local_pes_3_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_18_io_in_kv = local_pes_2_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_18_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_18_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_18_io_in_stage = local_pes_3_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_19_clock = clock;
  assign local_pes_3_19_reset = reset;
  assign local_pes_3_19_io_in_q = local_pes_3_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_19_io_in_sum = local_pes_3_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_19_io_in_sum_exp = local_pes_3_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_19_io_in_kv = local_pes_2_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_19_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_19_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_19_io_in_stage = local_pes_3_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_20_clock = clock;
  assign local_pes_3_20_reset = reset;
  assign local_pes_3_20_io_in_q = local_pes_3_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_20_io_in_sum = local_pes_3_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_20_io_in_sum_exp = local_pes_3_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_20_io_in_kv = local_pes_2_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_20_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_20_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_20_io_in_stage = local_pes_3_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_21_clock = clock;
  assign local_pes_3_21_reset = reset;
  assign local_pes_3_21_io_in_q = local_pes_3_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_21_io_in_sum = local_pes_3_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_21_io_in_sum_exp = local_pes_3_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_21_io_in_kv = local_pes_2_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_21_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_21_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_21_io_in_stage = local_pes_3_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_22_clock = clock;
  assign local_pes_3_22_reset = reset;
  assign local_pes_3_22_io_in_q = local_pes_3_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_22_io_in_sum = local_pes_3_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_22_io_in_sum_exp = local_pes_3_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_22_io_in_kv = local_pes_2_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_22_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_22_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_22_io_in_stage = local_pes_3_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_23_clock = clock;
  assign local_pes_3_23_reset = reset;
  assign local_pes_3_23_io_in_q = local_pes_3_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_23_io_in_sum = local_pes_3_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_23_io_in_sum_exp = local_pes_3_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_23_io_in_kv = local_pes_2_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_23_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_23_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_23_io_in_stage = local_pes_3_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_24_clock = clock;
  assign local_pes_3_24_reset = reset;
  assign local_pes_3_24_io_in_q = local_pes_3_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_24_io_in_sum = local_pes_3_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_24_io_in_sum_exp = local_pes_3_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_24_io_in_kv = local_pes_2_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_24_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_24_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_24_io_in_stage = local_pes_3_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_25_clock = clock;
  assign local_pes_3_25_reset = reset;
  assign local_pes_3_25_io_in_q = local_pes_3_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_25_io_in_sum = local_pes_3_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_25_io_in_sum_exp = local_pes_3_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_25_io_in_kv = local_pes_2_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_25_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_25_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_25_io_in_stage = local_pes_3_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_26_clock = clock;
  assign local_pes_3_26_reset = reset;
  assign local_pes_3_26_io_in_q = local_pes_3_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_26_io_in_sum = local_pes_3_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_26_io_in_sum_exp = local_pes_3_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_26_io_in_kv = local_pes_2_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_26_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_26_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_26_io_in_stage = local_pes_3_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_27_clock = clock;
  assign local_pes_3_27_reset = reset;
  assign local_pes_3_27_io_in_q = local_pes_3_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_27_io_in_sum = local_pes_3_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_27_io_in_sum_exp = local_pes_3_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_27_io_in_kv = local_pes_2_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_27_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_27_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_27_io_in_stage = local_pes_3_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_28_clock = clock;
  assign local_pes_3_28_reset = reset;
  assign local_pes_3_28_io_in_q = local_pes_3_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_28_io_in_sum = local_pes_3_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_28_io_in_sum_exp = local_pes_3_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_28_io_in_kv = local_pes_2_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_28_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_28_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_28_io_in_stage = local_pes_3_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_29_clock = clock;
  assign local_pes_3_29_reset = reset;
  assign local_pes_3_29_io_in_q = local_pes_3_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_29_io_in_sum = local_pes_3_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_29_io_in_sum_exp = local_pes_3_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_29_io_in_kv = local_pes_2_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_29_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_29_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_29_io_in_stage = local_pes_3_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_30_clock = clock;
  assign local_pes_3_30_reset = reset;
  assign local_pes_3_30_io_in_q = local_pes_3_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_30_io_in_sum = local_pes_3_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_30_io_in_sum_exp = local_pes_3_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_30_io_in_kv = local_pes_2_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_30_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_30_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_30_io_in_stage = local_pes_3_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_3_31_clock = clock;
  assign local_pes_3_31_reset = reset;
  assign local_pes_3_31_io_in_q = local_pes_3_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_3_31_io_in_sum = local_pes_3_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_3_31_io_in_sum_exp = local_pes_3_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_3_31_io_in_kv = local_pes_2_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_3_31_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_3_31_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_3_31_io_in_stage = local_pes_3_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_0_clock = clock;
  assign local_pes_4_0_reset = reset;
  assign local_pes_4_0_io_in_q = io_q_ports_4; // @[PEArray.scala 51:37]
  assign local_pes_4_0_io_in_kv = io_kv_ports_35; // @[PEArray.scala 40:34]
  assign local_pes_4_0_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_0_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_0_io_in_stage = io_stage_ports_4; // @[PEArray.scala 52:41]
  assign local_pes_4_1_clock = clock;
  assign local_pes_4_1_reset = reset;
  assign local_pes_4_1_io_in_q = local_pes_4_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_1_io_in_sum = local_pes_4_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_4_1_io_in_kv = local_pes_3_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_1_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_1_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_1_io_in_stage = local_pes_4_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_2_clock = clock;
  assign local_pes_4_2_reset = reset;
  assign local_pes_4_2_io_in_q = local_pes_4_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_2_io_in_sum = local_pes_4_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_2_io_in_sum_exp = local_pes_4_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_2_io_in_kv = local_pes_3_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_2_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_2_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_2_io_in_stage = local_pes_4_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_3_clock = clock;
  assign local_pes_4_3_reset = reset;
  assign local_pes_4_3_io_in_q = local_pes_4_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_3_io_in_sum = local_pes_4_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_3_io_in_sum_exp = local_pes_4_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_3_io_in_kv = local_pes_3_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_3_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_3_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_3_io_in_stage = local_pes_4_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_4_clock = clock;
  assign local_pes_4_4_reset = reset;
  assign local_pes_4_4_io_in_q = local_pes_4_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_4_io_in_sum = local_pes_4_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_4_io_in_sum_exp = local_pes_4_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_4_io_in_kv = local_pes_3_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_4_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_4_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_4_io_in_stage = local_pes_4_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_5_clock = clock;
  assign local_pes_4_5_reset = reset;
  assign local_pes_4_5_io_in_q = local_pes_4_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_5_io_in_sum = local_pes_4_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_5_io_in_sum_exp = local_pes_4_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_5_io_in_kv = local_pes_3_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_5_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_5_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_5_io_in_stage = local_pes_4_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_6_clock = clock;
  assign local_pes_4_6_reset = reset;
  assign local_pes_4_6_io_in_q = local_pes_4_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_6_io_in_sum = local_pes_4_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_6_io_in_sum_exp = local_pes_4_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_6_io_in_kv = local_pes_3_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_6_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_6_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_6_io_in_stage = local_pes_4_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_7_clock = clock;
  assign local_pes_4_7_reset = reset;
  assign local_pes_4_7_io_in_q = local_pes_4_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_7_io_in_sum = local_pes_4_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_7_io_in_sum_exp = local_pes_4_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_7_io_in_kv = local_pes_3_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_7_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_7_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_7_io_in_stage = local_pes_4_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_8_clock = clock;
  assign local_pes_4_8_reset = reset;
  assign local_pes_4_8_io_in_q = local_pes_4_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_8_io_in_sum = local_pes_4_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_8_io_in_sum_exp = local_pes_4_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_8_io_in_kv = local_pes_3_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_8_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_8_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_8_io_in_stage = local_pes_4_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_9_clock = clock;
  assign local_pes_4_9_reset = reset;
  assign local_pes_4_9_io_in_q = local_pes_4_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_9_io_in_sum = local_pes_4_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_9_io_in_sum_exp = local_pes_4_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_9_io_in_kv = local_pes_3_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_9_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_9_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_9_io_in_stage = local_pes_4_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_10_clock = clock;
  assign local_pes_4_10_reset = reset;
  assign local_pes_4_10_io_in_q = local_pes_4_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_10_io_in_sum = local_pes_4_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_10_io_in_sum_exp = local_pes_4_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_10_io_in_kv = local_pes_3_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_10_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_10_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_10_io_in_stage = local_pes_4_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_11_clock = clock;
  assign local_pes_4_11_reset = reset;
  assign local_pes_4_11_io_in_q = local_pes_4_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_11_io_in_sum = local_pes_4_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_11_io_in_sum_exp = local_pes_4_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_11_io_in_kv = local_pes_3_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_11_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_11_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_11_io_in_stage = local_pes_4_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_12_clock = clock;
  assign local_pes_4_12_reset = reset;
  assign local_pes_4_12_io_in_q = local_pes_4_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_12_io_in_sum = local_pes_4_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_12_io_in_sum_exp = local_pes_4_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_12_io_in_kv = local_pes_3_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_12_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_12_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_12_io_in_stage = local_pes_4_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_13_clock = clock;
  assign local_pes_4_13_reset = reset;
  assign local_pes_4_13_io_in_q = local_pes_4_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_13_io_in_sum = local_pes_4_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_13_io_in_sum_exp = local_pes_4_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_13_io_in_kv = local_pes_3_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_13_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_13_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_13_io_in_stage = local_pes_4_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_14_clock = clock;
  assign local_pes_4_14_reset = reset;
  assign local_pes_4_14_io_in_q = local_pes_4_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_14_io_in_sum = local_pes_4_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_14_io_in_sum_exp = local_pes_4_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_14_io_in_kv = local_pes_3_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_14_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_14_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_14_io_in_stage = local_pes_4_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_15_clock = clock;
  assign local_pes_4_15_reset = reset;
  assign local_pes_4_15_io_in_q = local_pes_4_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_15_io_in_sum = local_pes_4_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_15_io_in_sum_exp = local_pes_4_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_15_io_in_kv = local_pes_3_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_15_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_15_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_15_io_in_stage = local_pes_4_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_16_clock = clock;
  assign local_pes_4_16_reset = reset;
  assign local_pes_4_16_io_in_q = local_pes_4_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_16_io_in_sum = local_pes_4_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_16_io_in_sum_exp = local_pes_4_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_16_io_in_kv = local_pes_3_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_16_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_16_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_16_io_in_stage = local_pes_4_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_17_clock = clock;
  assign local_pes_4_17_reset = reset;
  assign local_pes_4_17_io_in_q = local_pes_4_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_17_io_in_sum = local_pes_4_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_17_io_in_sum_exp = local_pes_4_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_17_io_in_kv = local_pes_3_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_17_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_17_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_17_io_in_stage = local_pes_4_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_18_clock = clock;
  assign local_pes_4_18_reset = reset;
  assign local_pes_4_18_io_in_q = local_pes_4_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_18_io_in_sum = local_pes_4_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_18_io_in_sum_exp = local_pes_4_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_18_io_in_kv = local_pes_3_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_18_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_18_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_18_io_in_stage = local_pes_4_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_19_clock = clock;
  assign local_pes_4_19_reset = reset;
  assign local_pes_4_19_io_in_q = local_pes_4_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_19_io_in_sum = local_pes_4_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_19_io_in_sum_exp = local_pes_4_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_19_io_in_kv = local_pes_3_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_19_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_19_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_19_io_in_stage = local_pes_4_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_20_clock = clock;
  assign local_pes_4_20_reset = reset;
  assign local_pes_4_20_io_in_q = local_pes_4_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_20_io_in_sum = local_pes_4_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_20_io_in_sum_exp = local_pes_4_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_20_io_in_kv = local_pes_3_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_20_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_20_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_20_io_in_stage = local_pes_4_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_21_clock = clock;
  assign local_pes_4_21_reset = reset;
  assign local_pes_4_21_io_in_q = local_pes_4_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_21_io_in_sum = local_pes_4_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_21_io_in_sum_exp = local_pes_4_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_21_io_in_kv = local_pes_3_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_21_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_21_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_21_io_in_stage = local_pes_4_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_22_clock = clock;
  assign local_pes_4_22_reset = reset;
  assign local_pes_4_22_io_in_q = local_pes_4_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_22_io_in_sum = local_pes_4_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_22_io_in_sum_exp = local_pes_4_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_22_io_in_kv = local_pes_3_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_22_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_22_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_22_io_in_stage = local_pes_4_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_23_clock = clock;
  assign local_pes_4_23_reset = reset;
  assign local_pes_4_23_io_in_q = local_pes_4_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_23_io_in_sum = local_pes_4_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_23_io_in_sum_exp = local_pes_4_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_23_io_in_kv = local_pes_3_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_23_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_23_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_23_io_in_stage = local_pes_4_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_24_clock = clock;
  assign local_pes_4_24_reset = reset;
  assign local_pes_4_24_io_in_q = local_pes_4_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_24_io_in_sum = local_pes_4_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_24_io_in_sum_exp = local_pes_4_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_24_io_in_kv = local_pes_3_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_24_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_24_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_24_io_in_stage = local_pes_4_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_25_clock = clock;
  assign local_pes_4_25_reset = reset;
  assign local_pes_4_25_io_in_q = local_pes_4_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_25_io_in_sum = local_pes_4_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_25_io_in_sum_exp = local_pes_4_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_25_io_in_kv = local_pes_3_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_25_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_25_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_25_io_in_stage = local_pes_4_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_26_clock = clock;
  assign local_pes_4_26_reset = reset;
  assign local_pes_4_26_io_in_q = local_pes_4_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_26_io_in_sum = local_pes_4_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_26_io_in_sum_exp = local_pes_4_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_26_io_in_kv = local_pes_3_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_26_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_26_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_26_io_in_stage = local_pes_4_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_27_clock = clock;
  assign local_pes_4_27_reset = reset;
  assign local_pes_4_27_io_in_q = local_pes_4_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_27_io_in_sum = local_pes_4_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_27_io_in_sum_exp = local_pes_4_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_27_io_in_kv = local_pes_3_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_27_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_27_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_27_io_in_stage = local_pes_4_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_28_clock = clock;
  assign local_pes_4_28_reset = reset;
  assign local_pes_4_28_io_in_q = local_pes_4_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_28_io_in_sum = local_pes_4_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_28_io_in_sum_exp = local_pes_4_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_28_io_in_kv = local_pes_3_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_28_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_28_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_28_io_in_stage = local_pes_4_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_29_clock = clock;
  assign local_pes_4_29_reset = reset;
  assign local_pes_4_29_io_in_q = local_pes_4_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_29_io_in_sum = local_pes_4_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_29_io_in_sum_exp = local_pes_4_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_29_io_in_kv = local_pes_3_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_29_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_29_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_29_io_in_stage = local_pes_4_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_30_clock = clock;
  assign local_pes_4_30_reset = reset;
  assign local_pes_4_30_io_in_q = local_pes_4_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_30_io_in_sum = local_pes_4_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_30_io_in_sum_exp = local_pes_4_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_30_io_in_kv = local_pes_3_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_30_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_30_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_30_io_in_stage = local_pes_4_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_4_31_clock = clock;
  assign local_pes_4_31_reset = reset;
  assign local_pes_4_31_io_in_q = local_pes_4_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_4_31_io_in_sum = local_pes_4_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_4_31_io_in_sum_exp = local_pes_4_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_4_31_io_in_kv = local_pes_3_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_4_31_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_4_31_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_4_31_io_in_stage = local_pes_4_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_0_clock = clock;
  assign local_pes_5_0_reset = reset;
  assign local_pes_5_0_io_in_q = io_q_ports_5; // @[PEArray.scala 51:37]
  assign local_pes_5_0_io_in_kv = io_kv_ports_36; // @[PEArray.scala 40:34]
  assign local_pes_5_0_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_0_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_0_io_in_stage = io_stage_ports_5; // @[PEArray.scala 52:41]
  assign local_pes_5_1_clock = clock;
  assign local_pes_5_1_reset = reset;
  assign local_pes_5_1_io_in_q = local_pes_5_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_1_io_in_sum = local_pes_5_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_5_1_io_in_kv = local_pes_4_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_1_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_1_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_1_io_in_stage = local_pes_5_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_2_clock = clock;
  assign local_pes_5_2_reset = reset;
  assign local_pes_5_2_io_in_q = local_pes_5_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_2_io_in_sum = local_pes_5_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_2_io_in_sum_exp = local_pes_5_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_2_io_in_kv = local_pes_4_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_2_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_2_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_2_io_in_stage = local_pes_5_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_3_clock = clock;
  assign local_pes_5_3_reset = reset;
  assign local_pes_5_3_io_in_q = local_pes_5_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_3_io_in_sum = local_pes_5_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_3_io_in_sum_exp = local_pes_5_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_3_io_in_kv = local_pes_4_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_3_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_3_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_3_io_in_stage = local_pes_5_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_4_clock = clock;
  assign local_pes_5_4_reset = reset;
  assign local_pes_5_4_io_in_q = local_pes_5_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_4_io_in_sum = local_pes_5_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_4_io_in_sum_exp = local_pes_5_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_4_io_in_kv = local_pes_4_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_4_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_4_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_4_io_in_stage = local_pes_5_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_5_clock = clock;
  assign local_pes_5_5_reset = reset;
  assign local_pes_5_5_io_in_q = local_pes_5_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_5_io_in_sum = local_pes_5_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_5_io_in_sum_exp = local_pes_5_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_5_io_in_kv = local_pes_4_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_5_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_5_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_5_io_in_stage = local_pes_5_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_6_clock = clock;
  assign local_pes_5_6_reset = reset;
  assign local_pes_5_6_io_in_q = local_pes_5_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_6_io_in_sum = local_pes_5_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_6_io_in_sum_exp = local_pes_5_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_6_io_in_kv = local_pes_4_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_6_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_6_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_6_io_in_stage = local_pes_5_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_7_clock = clock;
  assign local_pes_5_7_reset = reset;
  assign local_pes_5_7_io_in_q = local_pes_5_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_7_io_in_sum = local_pes_5_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_7_io_in_sum_exp = local_pes_5_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_7_io_in_kv = local_pes_4_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_7_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_7_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_7_io_in_stage = local_pes_5_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_8_clock = clock;
  assign local_pes_5_8_reset = reset;
  assign local_pes_5_8_io_in_q = local_pes_5_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_8_io_in_sum = local_pes_5_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_8_io_in_sum_exp = local_pes_5_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_8_io_in_kv = local_pes_4_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_8_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_8_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_8_io_in_stage = local_pes_5_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_9_clock = clock;
  assign local_pes_5_9_reset = reset;
  assign local_pes_5_9_io_in_q = local_pes_5_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_9_io_in_sum = local_pes_5_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_9_io_in_sum_exp = local_pes_5_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_9_io_in_kv = local_pes_4_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_9_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_9_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_9_io_in_stage = local_pes_5_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_10_clock = clock;
  assign local_pes_5_10_reset = reset;
  assign local_pes_5_10_io_in_q = local_pes_5_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_10_io_in_sum = local_pes_5_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_10_io_in_sum_exp = local_pes_5_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_10_io_in_kv = local_pes_4_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_10_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_10_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_10_io_in_stage = local_pes_5_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_11_clock = clock;
  assign local_pes_5_11_reset = reset;
  assign local_pes_5_11_io_in_q = local_pes_5_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_11_io_in_sum = local_pes_5_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_11_io_in_sum_exp = local_pes_5_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_11_io_in_kv = local_pes_4_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_11_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_11_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_11_io_in_stage = local_pes_5_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_12_clock = clock;
  assign local_pes_5_12_reset = reset;
  assign local_pes_5_12_io_in_q = local_pes_5_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_12_io_in_sum = local_pes_5_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_12_io_in_sum_exp = local_pes_5_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_12_io_in_kv = local_pes_4_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_12_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_12_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_12_io_in_stage = local_pes_5_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_13_clock = clock;
  assign local_pes_5_13_reset = reset;
  assign local_pes_5_13_io_in_q = local_pes_5_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_13_io_in_sum = local_pes_5_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_13_io_in_sum_exp = local_pes_5_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_13_io_in_kv = local_pes_4_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_13_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_13_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_13_io_in_stage = local_pes_5_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_14_clock = clock;
  assign local_pes_5_14_reset = reset;
  assign local_pes_5_14_io_in_q = local_pes_5_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_14_io_in_sum = local_pes_5_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_14_io_in_sum_exp = local_pes_5_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_14_io_in_kv = local_pes_4_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_14_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_14_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_14_io_in_stage = local_pes_5_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_15_clock = clock;
  assign local_pes_5_15_reset = reset;
  assign local_pes_5_15_io_in_q = local_pes_5_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_15_io_in_sum = local_pes_5_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_15_io_in_sum_exp = local_pes_5_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_15_io_in_kv = local_pes_4_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_15_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_15_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_15_io_in_stage = local_pes_5_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_16_clock = clock;
  assign local_pes_5_16_reset = reset;
  assign local_pes_5_16_io_in_q = local_pes_5_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_16_io_in_sum = local_pes_5_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_16_io_in_sum_exp = local_pes_5_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_16_io_in_kv = local_pes_4_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_16_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_16_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_16_io_in_stage = local_pes_5_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_17_clock = clock;
  assign local_pes_5_17_reset = reset;
  assign local_pes_5_17_io_in_q = local_pes_5_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_17_io_in_sum = local_pes_5_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_17_io_in_sum_exp = local_pes_5_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_17_io_in_kv = local_pes_4_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_17_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_17_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_17_io_in_stage = local_pes_5_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_18_clock = clock;
  assign local_pes_5_18_reset = reset;
  assign local_pes_5_18_io_in_q = local_pes_5_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_18_io_in_sum = local_pes_5_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_18_io_in_sum_exp = local_pes_5_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_18_io_in_kv = local_pes_4_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_18_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_18_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_18_io_in_stage = local_pes_5_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_19_clock = clock;
  assign local_pes_5_19_reset = reset;
  assign local_pes_5_19_io_in_q = local_pes_5_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_19_io_in_sum = local_pes_5_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_19_io_in_sum_exp = local_pes_5_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_19_io_in_kv = local_pes_4_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_19_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_19_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_19_io_in_stage = local_pes_5_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_20_clock = clock;
  assign local_pes_5_20_reset = reset;
  assign local_pes_5_20_io_in_q = local_pes_5_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_20_io_in_sum = local_pes_5_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_20_io_in_sum_exp = local_pes_5_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_20_io_in_kv = local_pes_4_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_20_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_20_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_20_io_in_stage = local_pes_5_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_21_clock = clock;
  assign local_pes_5_21_reset = reset;
  assign local_pes_5_21_io_in_q = local_pes_5_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_21_io_in_sum = local_pes_5_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_21_io_in_sum_exp = local_pes_5_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_21_io_in_kv = local_pes_4_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_21_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_21_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_21_io_in_stage = local_pes_5_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_22_clock = clock;
  assign local_pes_5_22_reset = reset;
  assign local_pes_5_22_io_in_q = local_pes_5_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_22_io_in_sum = local_pes_5_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_22_io_in_sum_exp = local_pes_5_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_22_io_in_kv = local_pes_4_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_22_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_22_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_22_io_in_stage = local_pes_5_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_23_clock = clock;
  assign local_pes_5_23_reset = reset;
  assign local_pes_5_23_io_in_q = local_pes_5_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_23_io_in_sum = local_pes_5_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_23_io_in_sum_exp = local_pes_5_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_23_io_in_kv = local_pes_4_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_23_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_23_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_23_io_in_stage = local_pes_5_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_24_clock = clock;
  assign local_pes_5_24_reset = reset;
  assign local_pes_5_24_io_in_q = local_pes_5_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_24_io_in_sum = local_pes_5_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_24_io_in_sum_exp = local_pes_5_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_24_io_in_kv = local_pes_4_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_24_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_24_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_24_io_in_stage = local_pes_5_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_25_clock = clock;
  assign local_pes_5_25_reset = reset;
  assign local_pes_5_25_io_in_q = local_pes_5_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_25_io_in_sum = local_pes_5_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_25_io_in_sum_exp = local_pes_5_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_25_io_in_kv = local_pes_4_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_25_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_25_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_25_io_in_stage = local_pes_5_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_26_clock = clock;
  assign local_pes_5_26_reset = reset;
  assign local_pes_5_26_io_in_q = local_pes_5_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_26_io_in_sum = local_pes_5_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_26_io_in_sum_exp = local_pes_5_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_26_io_in_kv = local_pes_4_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_26_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_26_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_26_io_in_stage = local_pes_5_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_27_clock = clock;
  assign local_pes_5_27_reset = reset;
  assign local_pes_5_27_io_in_q = local_pes_5_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_27_io_in_sum = local_pes_5_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_27_io_in_sum_exp = local_pes_5_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_27_io_in_kv = local_pes_4_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_27_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_27_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_27_io_in_stage = local_pes_5_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_28_clock = clock;
  assign local_pes_5_28_reset = reset;
  assign local_pes_5_28_io_in_q = local_pes_5_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_28_io_in_sum = local_pes_5_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_28_io_in_sum_exp = local_pes_5_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_28_io_in_kv = local_pes_4_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_28_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_28_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_28_io_in_stage = local_pes_5_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_29_clock = clock;
  assign local_pes_5_29_reset = reset;
  assign local_pes_5_29_io_in_q = local_pes_5_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_29_io_in_sum = local_pes_5_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_29_io_in_sum_exp = local_pes_5_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_29_io_in_kv = local_pes_4_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_29_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_29_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_29_io_in_stage = local_pes_5_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_30_clock = clock;
  assign local_pes_5_30_reset = reset;
  assign local_pes_5_30_io_in_q = local_pes_5_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_30_io_in_sum = local_pes_5_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_30_io_in_sum_exp = local_pes_5_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_30_io_in_kv = local_pes_4_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_30_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_30_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_30_io_in_stage = local_pes_5_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_5_31_clock = clock;
  assign local_pes_5_31_reset = reset;
  assign local_pes_5_31_io_in_q = local_pes_5_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_5_31_io_in_sum = local_pes_5_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_5_31_io_in_sum_exp = local_pes_5_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_5_31_io_in_kv = local_pes_4_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_5_31_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_5_31_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_5_31_io_in_stage = local_pes_5_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_0_clock = clock;
  assign local_pes_6_0_reset = reset;
  assign local_pes_6_0_io_in_q = io_q_ports_6; // @[PEArray.scala 51:37]
  assign local_pes_6_0_io_in_kv = io_kv_ports_37; // @[PEArray.scala 40:34]
  assign local_pes_6_0_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_0_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_0_io_in_stage = io_stage_ports_6; // @[PEArray.scala 52:41]
  assign local_pes_6_1_clock = clock;
  assign local_pes_6_1_reset = reset;
  assign local_pes_6_1_io_in_q = local_pes_6_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_1_io_in_sum = local_pes_6_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_6_1_io_in_kv = local_pes_5_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_1_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_1_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_1_io_in_stage = local_pes_6_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_2_clock = clock;
  assign local_pes_6_2_reset = reset;
  assign local_pes_6_2_io_in_q = local_pes_6_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_2_io_in_sum = local_pes_6_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_2_io_in_sum_exp = local_pes_6_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_2_io_in_kv = local_pes_5_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_2_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_2_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_2_io_in_stage = local_pes_6_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_3_clock = clock;
  assign local_pes_6_3_reset = reset;
  assign local_pes_6_3_io_in_q = local_pes_6_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_3_io_in_sum = local_pes_6_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_3_io_in_sum_exp = local_pes_6_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_3_io_in_kv = local_pes_5_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_3_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_3_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_3_io_in_stage = local_pes_6_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_4_clock = clock;
  assign local_pes_6_4_reset = reset;
  assign local_pes_6_4_io_in_q = local_pes_6_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_4_io_in_sum = local_pes_6_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_4_io_in_sum_exp = local_pes_6_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_4_io_in_kv = local_pes_5_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_4_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_4_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_4_io_in_stage = local_pes_6_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_5_clock = clock;
  assign local_pes_6_5_reset = reset;
  assign local_pes_6_5_io_in_q = local_pes_6_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_5_io_in_sum = local_pes_6_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_5_io_in_sum_exp = local_pes_6_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_5_io_in_kv = local_pes_5_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_5_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_5_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_5_io_in_stage = local_pes_6_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_6_clock = clock;
  assign local_pes_6_6_reset = reset;
  assign local_pes_6_6_io_in_q = local_pes_6_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_6_io_in_sum = local_pes_6_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_6_io_in_sum_exp = local_pes_6_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_6_io_in_kv = local_pes_5_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_6_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_6_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_6_io_in_stage = local_pes_6_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_7_clock = clock;
  assign local_pes_6_7_reset = reset;
  assign local_pes_6_7_io_in_q = local_pes_6_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_7_io_in_sum = local_pes_6_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_7_io_in_sum_exp = local_pes_6_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_7_io_in_kv = local_pes_5_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_7_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_7_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_7_io_in_stage = local_pes_6_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_8_clock = clock;
  assign local_pes_6_8_reset = reset;
  assign local_pes_6_8_io_in_q = local_pes_6_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_8_io_in_sum = local_pes_6_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_8_io_in_sum_exp = local_pes_6_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_8_io_in_kv = local_pes_5_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_8_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_8_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_8_io_in_stage = local_pes_6_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_9_clock = clock;
  assign local_pes_6_9_reset = reset;
  assign local_pes_6_9_io_in_q = local_pes_6_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_9_io_in_sum = local_pes_6_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_9_io_in_sum_exp = local_pes_6_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_9_io_in_kv = local_pes_5_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_9_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_9_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_9_io_in_stage = local_pes_6_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_10_clock = clock;
  assign local_pes_6_10_reset = reset;
  assign local_pes_6_10_io_in_q = local_pes_6_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_10_io_in_sum = local_pes_6_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_10_io_in_sum_exp = local_pes_6_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_10_io_in_kv = local_pes_5_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_10_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_10_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_10_io_in_stage = local_pes_6_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_11_clock = clock;
  assign local_pes_6_11_reset = reset;
  assign local_pes_6_11_io_in_q = local_pes_6_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_11_io_in_sum = local_pes_6_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_11_io_in_sum_exp = local_pes_6_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_11_io_in_kv = local_pes_5_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_11_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_11_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_11_io_in_stage = local_pes_6_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_12_clock = clock;
  assign local_pes_6_12_reset = reset;
  assign local_pes_6_12_io_in_q = local_pes_6_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_12_io_in_sum = local_pes_6_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_12_io_in_sum_exp = local_pes_6_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_12_io_in_kv = local_pes_5_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_12_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_12_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_12_io_in_stage = local_pes_6_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_13_clock = clock;
  assign local_pes_6_13_reset = reset;
  assign local_pes_6_13_io_in_q = local_pes_6_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_13_io_in_sum = local_pes_6_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_13_io_in_sum_exp = local_pes_6_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_13_io_in_kv = local_pes_5_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_13_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_13_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_13_io_in_stage = local_pes_6_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_14_clock = clock;
  assign local_pes_6_14_reset = reset;
  assign local_pes_6_14_io_in_q = local_pes_6_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_14_io_in_sum = local_pes_6_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_14_io_in_sum_exp = local_pes_6_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_14_io_in_kv = local_pes_5_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_14_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_14_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_14_io_in_stage = local_pes_6_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_15_clock = clock;
  assign local_pes_6_15_reset = reset;
  assign local_pes_6_15_io_in_q = local_pes_6_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_15_io_in_sum = local_pes_6_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_15_io_in_sum_exp = local_pes_6_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_15_io_in_kv = local_pes_5_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_15_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_15_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_15_io_in_stage = local_pes_6_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_16_clock = clock;
  assign local_pes_6_16_reset = reset;
  assign local_pes_6_16_io_in_q = local_pes_6_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_16_io_in_sum = local_pes_6_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_16_io_in_sum_exp = local_pes_6_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_16_io_in_kv = local_pes_5_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_16_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_16_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_16_io_in_stage = local_pes_6_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_17_clock = clock;
  assign local_pes_6_17_reset = reset;
  assign local_pes_6_17_io_in_q = local_pes_6_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_17_io_in_sum = local_pes_6_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_17_io_in_sum_exp = local_pes_6_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_17_io_in_kv = local_pes_5_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_17_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_17_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_17_io_in_stage = local_pes_6_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_18_clock = clock;
  assign local_pes_6_18_reset = reset;
  assign local_pes_6_18_io_in_q = local_pes_6_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_18_io_in_sum = local_pes_6_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_18_io_in_sum_exp = local_pes_6_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_18_io_in_kv = local_pes_5_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_18_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_18_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_18_io_in_stage = local_pes_6_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_19_clock = clock;
  assign local_pes_6_19_reset = reset;
  assign local_pes_6_19_io_in_q = local_pes_6_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_19_io_in_sum = local_pes_6_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_19_io_in_sum_exp = local_pes_6_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_19_io_in_kv = local_pes_5_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_19_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_19_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_19_io_in_stage = local_pes_6_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_20_clock = clock;
  assign local_pes_6_20_reset = reset;
  assign local_pes_6_20_io_in_q = local_pes_6_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_20_io_in_sum = local_pes_6_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_20_io_in_sum_exp = local_pes_6_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_20_io_in_kv = local_pes_5_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_20_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_20_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_20_io_in_stage = local_pes_6_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_21_clock = clock;
  assign local_pes_6_21_reset = reset;
  assign local_pes_6_21_io_in_q = local_pes_6_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_21_io_in_sum = local_pes_6_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_21_io_in_sum_exp = local_pes_6_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_21_io_in_kv = local_pes_5_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_21_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_21_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_21_io_in_stage = local_pes_6_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_22_clock = clock;
  assign local_pes_6_22_reset = reset;
  assign local_pes_6_22_io_in_q = local_pes_6_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_22_io_in_sum = local_pes_6_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_22_io_in_sum_exp = local_pes_6_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_22_io_in_kv = local_pes_5_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_22_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_22_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_22_io_in_stage = local_pes_6_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_23_clock = clock;
  assign local_pes_6_23_reset = reset;
  assign local_pes_6_23_io_in_q = local_pes_6_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_23_io_in_sum = local_pes_6_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_23_io_in_sum_exp = local_pes_6_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_23_io_in_kv = local_pes_5_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_23_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_23_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_23_io_in_stage = local_pes_6_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_24_clock = clock;
  assign local_pes_6_24_reset = reset;
  assign local_pes_6_24_io_in_q = local_pes_6_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_24_io_in_sum = local_pes_6_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_24_io_in_sum_exp = local_pes_6_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_24_io_in_kv = local_pes_5_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_24_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_24_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_24_io_in_stage = local_pes_6_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_25_clock = clock;
  assign local_pes_6_25_reset = reset;
  assign local_pes_6_25_io_in_q = local_pes_6_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_25_io_in_sum = local_pes_6_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_25_io_in_sum_exp = local_pes_6_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_25_io_in_kv = local_pes_5_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_25_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_25_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_25_io_in_stage = local_pes_6_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_26_clock = clock;
  assign local_pes_6_26_reset = reset;
  assign local_pes_6_26_io_in_q = local_pes_6_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_26_io_in_sum = local_pes_6_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_26_io_in_sum_exp = local_pes_6_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_26_io_in_kv = local_pes_5_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_26_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_26_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_26_io_in_stage = local_pes_6_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_27_clock = clock;
  assign local_pes_6_27_reset = reset;
  assign local_pes_6_27_io_in_q = local_pes_6_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_27_io_in_sum = local_pes_6_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_27_io_in_sum_exp = local_pes_6_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_27_io_in_kv = local_pes_5_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_27_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_27_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_27_io_in_stage = local_pes_6_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_28_clock = clock;
  assign local_pes_6_28_reset = reset;
  assign local_pes_6_28_io_in_q = local_pes_6_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_28_io_in_sum = local_pes_6_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_28_io_in_sum_exp = local_pes_6_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_28_io_in_kv = local_pes_5_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_28_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_28_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_28_io_in_stage = local_pes_6_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_29_clock = clock;
  assign local_pes_6_29_reset = reset;
  assign local_pes_6_29_io_in_q = local_pes_6_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_29_io_in_sum = local_pes_6_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_29_io_in_sum_exp = local_pes_6_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_29_io_in_kv = local_pes_5_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_29_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_29_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_29_io_in_stage = local_pes_6_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_30_clock = clock;
  assign local_pes_6_30_reset = reset;
  assign local_pes_6_30_io_in_q = local_pes_6_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_30_io_in_sum = local_pes_6_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_30_io_in_sum_exp = local_pes_6_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_30_io_in_kv = local_pes_5_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_30_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_30_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_30_io_in_stage = local_pes_6_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_6_31_clock = clock;
  assign local_pes_6_31_reset = reset;
  assign local_pes_6_31_io_in_q = local_pes_6_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_6_31_io_in_sum = local_pes_6_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_6_31_io_in_sum_exp = local_pes_6_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_6_31_io_in_kv = local_pes_5_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_6_31_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_6_31_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_6_31_io_in_stage = local_pes_6_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_0_clock = clock;
  assign local_pes_7_0_reset = reset;
  assign local_pes_7_0_io_in_q = io_q_ports_7; // @[PEArray.scala 51:37]
  assign local_pes_7_0_io_in_kv = io_kv_ports_38; // @[PEArray.scala 40:34]
  assign local_pes_7_0_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_0_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_0_io_in_stage = io_stage_ports_7; // @[PEArray.scala 52:41]
  assign local_pes_7_1_clock = clock;
  assign local_pes_7_1_reset = reset;
  assign local_pes_7_1_io_in_q = local_pes_7_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_1_io_in_sum = local_pes_7_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_7_1_io_in_kv = local_pes_6_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_1_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_1_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_1_io_in_stage = local_pes_7_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_2_clock = clock;
  assign local_pes_7_2_reset = reset;
  assign local_pes_7_2_io_in_q = local_pes_7_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_2_io_in_sum = local_pes_7_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_2_io_in_sum_exp = local_pes_7_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_2_io_in_kv = local_pes_6_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_2_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_2_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_2_io_in_stage = local_pes_7_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_3_clock = clock;
  assign local_pes_7_3_reset = reset;
  assign local_pes_7_3_io_in_q = local_pes_7_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_3_io_in_sum = local_pes_7_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_3_io_in_sum_exp = local_pes_7_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_3_io_in_kv = local_pes_6_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_3_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_3_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_3_io_in_stage = local_pes_7_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_4_clock = clock;
  assign local_pes_7_4_reset = reset;
  assign local_pes_7_4_io_in_q = local_pes_7_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_4_io_in_sum = local_pes_7_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_4_io_in_sum_exp = local_pes_7_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_4_io_in_kv = local_pes_6_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_4_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_4_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_4_io_in_stage = local_pes_7_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_5_clock = clock;
  assign local_pes_7_5_reset = reset;
  assign local_pes_7_5_io_in_q = local_pes_7_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_5_io_in_sum = local_pes_7_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_5_io_in_sum_exp = local_pes_7_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_5_io_in_kv = local_pes_6_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_5_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_5_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_5_io_in_stage = local_pes_7_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_6_clock = clock;
  assign local_pes_7_6_reset = reset;
  assign local_pes_7_6_io_in_q = local_pes_7_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_6_io_in_sum = local_pes_7_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_6_io_in_sum_exp = local_pes_7_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_6_io_in_kv = local_pes_6_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_6_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_6_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_6_io_in_stage = local_pes_7_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_7_clock = clock;
  assign local_pes_7_7_reset = reset;
  assign local_pes_7_7_io_in_q = local_pes_7_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_7_io_in_sum = local_pes_7_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_7_io_in_sum_exp = local_pes_7_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_7_io_in_kv = local_pes_6_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_7_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_7_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_7_io_in_stage = local_pes_7_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_8_clock = clock;
  assign local_pes_7_8_reset = reset;
  assign local_pes_7_8_io_in_q = local_pes_7_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_8_io_in_sum = local_pes_7_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_8_io_in_sum_exp = local_pes_7_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_8_io_in_kv = local_pes_6_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_8_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_8_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_8_io_in_stage = local_pes_7_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_9_clock = clock;
  assign local_pes_7_9_reset = reset;
  assign local_pes_7_9_io_in_q = local_pes_7_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_9_io_in_sum = local_pes_7_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_9_io_in_sum_exp = local_pes_7_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_9_io_in_kv = local_pes_6_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_9_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_9_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_9_io_in_stage = local_pes_7_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_10_clock = clock;
  assign local_pes_7_10_reset = reset;
  assign local_pes_7_10_io_in_q = local_pes_7_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_10_io_in_sum = local_pes_7_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_10_io_in_sum_exp = local_pes_7_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_10_io_in_kv = local_pes_6_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_10_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_10_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_10_io_in_stage = local_pes_7_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_11_clock = clock;
  assign local_pes_7_11_reset = reset;
  assign local_pes_7_11_io_in_q = local_pes_7_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_11_io_in_sum = local_pes_7_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_11_io_in_sum_exp = local_pes_7_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_11_io_in_kv = local_pes_6_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_11_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_11_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_11_io_in_stage = local_pes_7_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_12_clock = clock;
  assign local_pes_7_12_reset = reset;
  assign local_pes_7_12_io_in_q = local_pes_7_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_12_io_in_sum = local_pes_7_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_12_io_in_sum_exp = local_pes_7_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_12_io_in_kv = local_pes_6_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_12_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_12_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_12_io_in_stage = local_pes_7_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_13_clock = clock;
  assign local_pes_7_13_reset = reset;
  assign local_pes_7_13_io_in_q = local_pes_7_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_13_io_in_sum = local_pes_7_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_13_io_in_sum_exp = local_pes_7_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_13_io_in_kv = local_pes_6_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_13_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_13_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_13_io_in_stage = local_pes_7_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_14_clock = clock;
  assign local_pes_7_14_reset = reset;
  assign local_pes_7_14_io_in_q = local_pes_7_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_14_io_in_sum = local_pes_7_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_14_io_in_sum_exp = local_pes_7_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_14_io_in_kv = local_pes_6_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_14_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_14_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_14_io_in_stage = local_pes_7_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_15_clock = clock;
  assign local_pes_7_15_reset = reset;
  assign local_pes_7_15_io_in_q = local_pes_7_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_15_io_in_sum = local_pes_7_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_15_io_in_sum_exp = local_pes_7_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_15_io_in_kv = local_pes_6_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_15_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_15_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_15_io_in_stage = local_pes_7_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_16_clock = clock;
  assign local_pes_7_16_reset = reset;
  assign local_pes_7_16_io_in_q = local_pes_7_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_16_io_in_sum = local_pes_7_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_16_io_in_sum_exp = local_pes_7_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_16_io_in_kv = local_pes_6_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_16_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_16_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_16_io_in_stage = local_pes_7_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_17_clock = clock;
  assign local_pes_7_17_reset = reset;
  assign local_pes_7_17_io_in_q = local_pes_7_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_17_io_in_sum = local_pes_7_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_17_io_in_sum_exp = local_pes_7_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_17_io_in_kv = local_pes_6_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_17_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_17_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_17_io_in_stage = local_pes_7_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_18_clock = clock;
  assign local_pes_7_18_reset = reset;
  assign local_pes_7_18_io_in_q = local_pes_7_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_18_io_in_sum = local_pes_7_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_18_io_in_sum_exp = local_pes_7_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_18_io_in_kv = local_pes_6_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_18_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_18_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_18_io_in_stage = local_pes_7_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_19_clock = clock;
  assign local_pes_7_19_reset = reset;
  assign local_pes_7_19_io_in_q = local_pes_7_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_19_io_in_sum = local_pes_7_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_19_io_in_sum_exp = local_pes_7_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_19_io_in_kv = local_pes_6_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_19_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_19_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_19_io_in_stage = local_pes_7_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_20_clock = clock;
  assign local_pes_7_20_reset = reset;
  assign local_pes_7_20_io_in_q = local_pes_7_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_20_io_in_sum = local_pes_7_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_20_io_in_sum_exp = local_pes_7_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_20_io_in_kv = local_pes_6_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_20_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_20_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_20_io_in_stage = local_pes_7_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_21_clock = clock;
  assign local_pes_7_21_reset = reset;
  assign local_pes_7_21_io_in_q = local_pes_7_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_21_io_in_sum = local_pes_7_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_21_io_in_sum_exp = local_pes_7_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_21_io_in_kv = local_pes_6_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_21_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_21_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_21_io_in_stage = local_pes_7_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_22_clock = clock;
  assign local_pes_7_22_reset = reset;
  assign local_pes_7_22_io_in_q = local_pes_7_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_22_io_in_sum = local_pes_7_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_22_io_in_sum_exp = local_pes_7_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_22_io_in_kv = local_pes_6_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_22_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_22_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_22_io_in_stage = local_pes_7_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_23_clock = clock;
  assign local_pes_7_23_reset = reset;
  assign local_pes_7_23_io_in_q = local_pes_7_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_23_io_in_sum = local_pes_7_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_23_io_in_sum_exp = local_pes_7_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_23_io_in_kv = local_pes_6_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_23_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_23_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_23_io_in_stage = local_pes_7_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_24_clock = clock;
  assign local_pes_7_24_reset = reset;
  assign local_pes_7_24_io_in_q = local_pes_7_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_24_io_in_sum = local_pes_7_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_24_io_in_sum_exp = local_pes_7_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_24_io_in_kv = local_pes_6_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_24_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_24_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_24_io_in_stage = local_pes_7_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_25_clock = clock;
  assign local_pes_7_25_reset = reset;
  assign local_pes_7_25_io_in_q = local_pes_7_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_25_io_in_sum = local_pes_7_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_25_io_in_sum_exp = local_pes_7_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_25_io_in_kv = local_pes_6_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_25_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_25_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_25_io_in_stage = local_pes_7_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_26_clock = clock;
  assign local_pes_7_26_reset = reset;
  assign local_pes_7_26_io_in_q = local_pes_7_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_26_io_in_sum = local_pes_7_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_26_io_in_sum_exp = local_pes_7_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_26_io_in_kv = local_pes_6_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_26_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_26_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_26_io_in_stage = local_pes_7_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_27_clock = clock;
  assign local_pes_7_27_reset = reset;
  assign local_pes_7_27_io_in_q = local_pes_7_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_27_io_in_sum = local_pes_7_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_27_io_in_sum_exp = local_pes_7_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_27_io_in_kv = local_pes_6_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_27_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_27_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_27_io_in_stage = local_pes_7_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_28_clock = clock;
  assign local_pes_7_28_reset = reset;
  assign local_pes_7_28_io_in_q = local_pes_7_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_28_io_in_sum = local_pes_7_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_28_io_in_sum_exp = local_pes_7_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_28_io_in_kv = local_pes_6_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_28_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_28_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_28_io_in_stage = local_pes_7_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_29_clock = clock;
  assign local_pes_7_29_reset = reset;
  assign local_pes_7_29_io_in_q = local_pes_7_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_29_io_in_sum = local_pes_7_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_29_io_in_sum_exp = local_pes_7_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_29_io_in_kv = local_pes_6_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_29_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_29_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_29_io_in_stage = local_pes_7_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_30_clock = clock;
  assign local_pes_7_30_reset = reset;
  assign local_pes_7_30_io_in_q = local_pes_7_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_30_io_in_sum = local_pes_7_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_30_io_in_sum_exp = local_pes_7_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_30_io_in_kv = local_pes_6_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_30_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_30_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_30_io_in_stage = local_pes_7_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_7_31_clock = clock;
  assign local_pes_7_31_reset = reset;
  assign local_pes_7_31_io_in_q = local_pes_7_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_7_31_io_in_sum = local_pes_7_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_7_31_io_in_sum_exp = local_pes_7_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_7_31_io_in_kv = local_pes_6_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_7_31_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_7_31_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_7_31_io_in_stage = local_pes_7_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_0_clock = clock;
  assign local_pes_8_0_reset = reset;
  assign local_pes_8_0_io_in_q = io_q_ports_8; // @[PEArray.scala 51:37]
  assign local_pes_8_0_io_in_kv = io_kv_ports_39; // @[PEArray.scala 40:34]
  assign local_pes_8_0_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_0_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_0_io_in_stage = io_stage_ports_8; // @[PEArray.scala 52:41]
  assign local_pes_8_1_clock = clock;
  assign local_pes_8_1_reset = reset;
  assign local_pes_8_1_io_in_q = local_pes_8_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_1_io_in_sum = local_pes_8_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_8_1_io_in_kv = local_pes_7_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_1_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_1_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_1_io_in_stage = local_pes_8_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_2_clock = clock;
  assign local_pes_8_2_reset = reset;
  assign local_pes_8_2_io_in_q = local_pes_8_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_2_io_in_sum = local_pes_8_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_2_io_in_sum_exp = local_pes_8_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_2_io_in_kv = local_pes_7_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_2_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_2_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_2_io_in_stage = local_pes_8_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_3_clock = clock;
  assign local_pes_8_3_reset = reset;
  assign local_pes_8_3_io_in_q = local_pes_8_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_3_io_in_sum = local_pes_8_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_3_io_in_sum_exp = local_pes_8_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_3_io_in_kv = local_pes_7_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_3_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_3_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_3_io_in_stage = local_pes_8_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_4_clock = clock;
  assign local_pes_8_4_reset = reset;
  assign local_pes_8_4_io_in_q = local_pes_8_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_4_io_in_sum = local_pes_8_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_4_io_in_sum_exp = local_pes_8_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_4_io_in_kv = local_pes_7_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_4_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_4_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_4_io_in_stage = local_pes_8_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_5_clock = clock;
  assign local_pes_8_5_reset = reset;
  assign local_pes_8_5_io_in_q = local_pes_8_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_5_io_in_sum = local_pes_8_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_5_io_in_sum_exp = local_pes_8_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_5_io_in_kv = local_pes_7_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_5_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_5_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_5_io_in_stage = local_pes_8_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_6_clock = clock;
  assign local_pes_8_6_reset = reset;
  assign local_pes_8_6_io_in_q = local_pes_8_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_6_io_in_sum = local_pes_8_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_6_io_in_sum_exp = local_pes_8_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_6_io_in_kv = local_pes_7_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_6_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_6_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_6_io_in_stage = local_pes_8_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_7_clock = clock;
  assign local_pes_8_7_reset = reset;
  assign local_pes_8_7_io_in_q = local_pes_8_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_7_io_in_sum = local_pes_8_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_7_io_in_sum_exp = local_pes_8_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_7_io_in_kv = local_pes_7_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_7_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_7_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_7_io_in_stage = local_pes_8_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_8_clock = clock;
  assign local_pes_8_8_reset = reset;
  assign local_pes_8_8_io_in_q = local_pes_8_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_8_io_in_sum = local_pes_8_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_8_io_in_sum_exp = local_pes_8_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_8_io_in_kv = local_pes_7_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_8_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_8_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_8_io_in_stage = local_pes_8_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_9_clock = clock;
  assign local_pes_8_9_reset = reset;
  assign local_pes_8_9_io_in_q = local_pes_8_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_9_io_in_sum = local_pes_8_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_9_io_in_sum_exp = local_pes_8_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_9_io_in_kv = local_pes_7_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_9_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_9_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_9_io_in_stage = local_pes_8_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_10_clock = clock;
  assign local_pes_8_10_reset = reset;
  assign local_pes_8_10_io_in_q = local_pes_8_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_10_io_in_sum = local_pes_8_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_10_io_in_sum_exp = local_pes_8_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_10_io_in_kv = local_pes_7_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_10_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_10_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_10_io_in_stage = local_pes_8_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_11_clock = clock;
  assign local_pes_8_11_reset = reset;
  assign local_pes_8_11_io_in_q = local_pes_8_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_11_io_in_sum = local_pes_8_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_11_io_in_sum_exp = local_pes_8_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_11_io_in_kv = local_pes_7_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_11_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_11_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_11_io_in_stage = local_pes_8_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_12_clock = clock;
  assign local_pes_8_12_reset = reset;
  assign local_pes_8_12_io_in_q = local_pes_8_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_12_io_in_sum = local_pes_8_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_12_io_in_sum_exp = local_pes_8_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_12_io_in_kv = local_pes_7_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_12_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_12_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_12_io_in_stage = local_pes_8_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_13_clock = clock;
  assign local_pes_8_13_reset = reset;
  assign local_pes_8_13_io_in_q = local_pes_8_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_13_io_in_sum = local_pes_8_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_13_io_in_sum_exp = local_pes_8_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_13_io_in_kv = local_pes_7_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_13_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_13_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_13_io_in_stage = local_pes_8_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_14_clock = clock;
  assign local_pes_8_14_reset = reset;
  assign local_pes_8_14_io_in_q = local_pes_8_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_14_io_in_sum = local_pes_8_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_14_io_in_sum_exp = local_pes_8_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_14_io_in_kv = local_pes_7_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_14_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_14_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_14_io_in_stage = local_pes_8_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_15_clock = clock;
  assign local_pes_8_15_reset = reset;
  assign local_pes_8_15_io_in_q = local_pes_8_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_15_io_in_sum = local_pes_8_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_15_io_in_sum_exp = local_pes_8_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_15_io_in_kv = local_pes_7_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_15_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_15_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_15_io_in_stage = local_pes_8_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_16_clock = clock;
  assign local_pes_8_16_reset = reset;
  assign local_pes_8_16_io_in_q = local_pes_8_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_16_io_in_sum = local_pes_8_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_16_io_in_sum_exp = local_pes_8_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_16_io_in_kv = local_pes_7_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_16_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_16_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_16_io_in_stage = local_pes_8_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_17_clock = clock;
  assign local_pes_8_17_reset = reset;
  assign local_pes_8_17_io_in_q = local_pes_8_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_17_io_in_sum = local_pes_8_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_17_io_in_sum_exp = local_pes_8_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_17_io_in_kv = local_pes_7_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_17_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_17_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_17_io_in_stage = local_pes_8_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_18_clock = clock;
  assign local_pes_8_18_reset = reset;
  assign local_pes_8_18_io_in_q = local_pes_8_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_18_io_in_sum = local_pes_8_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_18_io_in_sum_exp = local_pes_8_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_18_io_in_kv = local_pes_7_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_18_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_18_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_18_io_in_stage = local_pes_8_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_19_clock = clock;
  assign local_pes_8_19_reset = reset;
  assign local_pes_8_19_io_in_q = local_pes_8_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_19_io_in_sum = local_pes_8_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_19_io_in_sum_exp = local_pes_8_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_19_io_in_kv = local_pes_7_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_19_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_19_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_19_io_in_stage = local_pes_8_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_20_clock = clock;
  assign local_pes_8_20_reset = reset;
  assign local_pes_8_20_io_in_q = local_pes_8_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_20_io_in_sum = local_pes_8_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_20_io_in_sum_exp = local_pes_8_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_20_io_in_kv = local_pes_7_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_20_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_20_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_20_io_in_stage = local_pes_8_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_21_clock = clock;
  assign local_pes_8_21_reset = reset;
  assign local_pes_8_21_io_in_q = local_pes_8_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_21_io_in_sum = local_pes_8_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_21_io_in_sum_exp = local_pes_8_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_21_io_in_kv = local_pes_7_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_21_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_21_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_21_io_in_stage = local_pes_8_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_22_clock = clock;
  assign local_pes_8_22_reset = reset;
  assign local_pes_8_22_io_in_q = local_pes_8_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_22_io_in_sum = local_pes_8_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_22_io_in_sum_exp = local_pes_8_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_22_io_in_kv = local_pes_7_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_22_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_22_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_22_io_in_stage = local_pes_8_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_23_clock = clock;
  assign local_pes_8_23_reset = reset;
  assign local_pes_8_23_io_in_q = local_pes_8_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_23_io_in_sum = local_pes_8_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_23_io_in_sum_exp = local_pes_8_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_23_io_in_kv = local_pes_7_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_23_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_23_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_23_io_in_stage = local_pes_8_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_24_clock = clock;
  assign local_pes_8_24_reset = reset;
  assign local_pes_8_24_io_in_q = local_pes_8_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_24_io_in_sum = local_pes_8_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_24_io_in_sum_exp = local_pes_8_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_24_io_in_kv = local_pes_7_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_24_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_24_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_24_io_in_stage = local_pes_8_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_25_clock = clock;
  assign local_pes_8_25_reset = reset;
  assign local_pes_8_25_io_in_q = local_pes_8_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_25_io_in_sum = local_pes_8_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_25_io_in_sum_exp = local_pes_8_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_25_io_in_kv = local_pes_7_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_25_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_25_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_25_io_in_stage = local_pes_8_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_26_clock = clock;
  assign local_pes_8_26_reset = reset;
  assign local_pes_8_26_io_in_q = local_pes_8_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_26_io_in_sum = local_pes_8_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_26_io_in_sum_exp = local_pes_8_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_26_io_in_kv = local_pes_7_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_26_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_26_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_26_io_in_stage = local_pes_8_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_27_clock = clock;
  assign local_pes_8_27_reset = reset;
  assign local_pes_8_27_io_in_q = local_pes_8_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_27_io_in_sum = local_pes_8_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_27_io_in_sum_exp = local_pes_8_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_27_io_in_kv = local_pes_7_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_27_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_27_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_27_io_in_stage = local_pes_8_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_28_clock = clock;
  assign local_pes_8_28_reset = reset;
  assign local_pes_8_28_io_in_q = local_pes_8_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_28_io_in_sum = local_pes_8_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_28_io_in_sum_exp = local_pes_8_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_28_io_in_kv = local_pes_7_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_28_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_28_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_28_io_in_stage = local_pes_8_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_29_clock = clock;
  assign local_pes_8_29_reset = reset;
  assign local_pes_8_29_io_in_q = local_pes_8_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_29_io_in_sum = local_pes_8_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_29_io_in_sum_exp = local_pes_8_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_29_io_in_kv = local_pes_7_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_29_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_29_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_29_io_in_stage = local_pes_8_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_30_clock = clock;
  assign local_pes_8_30_reset = reset;
  assign local_pes_8_30_io_in_q = local_pes_8_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_30_io_in_sum = local_pes_8_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_30_io_in_sum_exp = local_pes_8_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_30_io_in_kv = local_pes_7_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_30_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_30_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_30_io_in_stage = local_pes_8_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_8_31_clock = clock;
  assign local_pes_8_31_reset = reset;
  assign local_pes_8_31_io_in_q = local_pes_8_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_8_31_io_in_sum = local_pes_8_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_8_31_io_in_sum_exp = local_pes_8_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_8_31_io_in_kv = local_pes_7_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_8_31_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_8_31_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_8_31_io_in_stage = local_pes_8_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_0_clock = clock;
  assign local_pes_9_0_reset = reset;
  assign local_pes_9_0_io_in_q = io_q_ports_9; // @[PEArray.scala 51:37]
  assign local_pes_9_0_io_in_kv = io_kv_ports_40; // @[PEArray.scala 40:34]
  assign local_pes_9_0_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_0_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_0_io_in_stage = io_stage_ports_9; // @[PEArray.scala 52:41]
  assign local_pes_9_1_clock = clock;
  assign local_pes_9_1_reset = reset;
  assign local_pes_9_1_io_in_q = local_pes_9_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_1_io_in_sum = local_pes_9_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_9_1_io_in_kv = local_pes_8_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_1_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_1_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_1_io_in_stage = local_pes_9_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_2_clock = clock;
  assign local_pes_9_2_reset = reset;
  assign local_pes_9_2_io_in_q = local_pes_9_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_2_io_in_sum = local_pes_9_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_2_io_in_sum_exp = local_pes_9_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_2_io_in_kv = local_pes_8_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_2_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_2_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_2_io_in_stage = local_pes_9_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_3_clock = clock;
  assign local_pes_9_3_reset = reset;
  assign local_pes_9_3_io_in_q = local_pes_9_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_3_io_in_sum = local_pes_9_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_3_io_in_sum_exp = local_pes_9_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_3_io_in_kv = local_pes_8_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_3_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_3_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_3_io_in_stage = local_pes_9_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_4_clock = clock;
  assign local_pes_9_4_reset = reset;
  assign local_pes_9_4_io_in_q = local_pes_9_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_4_io_in_sum = local_pes_9_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_4_io_in_sum_exp = local_pes_9_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_4_io_in_kv = local_pes_8_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_4_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_4_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_4_io_in_stage = local_pes_9_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_5_clock = clock;
  assign local_pes_9_5_reset = reset;
  assign local_pes_9_5_io_in_q = local_pes_9_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_5_io_in_sum = local_pes_9_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_5_io_in_sum_exp = local_pes_9_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_5_io_in_kv = local_pes_8_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_5_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_5_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_5_io_in_stage = local_pes_9_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_6_clock = clock;
  assign local_pes_9_6_reset = reset;
  assign local_pes_9_6_io_in_q = local_pes_9_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_6_io_in_sum = local_pes_9_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_6_io_in_sum_exp = local_pes_9_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_6_io_in_kv = local_pes_8_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_6_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_6_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_6_io_in_stage = local_pes_9_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_7_clock = clock;
  assign local_pes_9_7_reset = reset;
  assign local_pes_9_7_io_in_q = local_pes_9_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_7_io_in_sum = local_pes_9_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_7_io_in_sum_exp = local_pes_9_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_7_io_in_kv = local_pes_8_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_7_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_7_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_7_io_in_stage = local_pes_9_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_8_clock = clock;
  assign local_pes_9_8_reset = reset;
  assign local_pes_9_8_io_in_q = local_pes_9_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_8_io_in_sum = local_pes_9_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_8_io_in_sum_exp = local_pes_9_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_8_io_in_kv = local_pes_8_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_8_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_8_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_8_io_in_stage = local_pes_9_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_9_clock = clock;
  assign local_pes_9_9_reset = reset;
  assign local_pes_9_9_io_in_q = local_pes_9_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_9_io_in_sum = local_pes_9_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_9_io_in_sum_exp = local_pes_9_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_9_io_in_kv = local_pes_8_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_9_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_9_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_9_io_in_stage = local_pes_9_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_10_clock = clock;
  assign local_pes_9_10_reset = reset;
  assign local_pes_9_10_io_in_q = local_pes_9_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_10_io_in_sum = local_pes_9_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_10_io_in_sum_exp = local_pes_9_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_10_io_in_kv = local_pes_8_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_10_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_10_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_10_io_in_stage = local_pes_9_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_11_clock = clock;
  assign local_pes_9_11_reset = reset;
  assign local_pes_9_11_io_in_q = local_pes_9_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_11_io_in_sum = local_pes_9_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_11_io_in_sum_exp = local_pes_9_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_11_io_in_kv = local_pes_8_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_11_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_11_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_11_io_in_stage = local_pes_9_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_12_clock = clock;
  assign local_pes_9_12_reset = reset;
  assign local_pes_9_12_io_in_q = local_pes_9_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_12_io_in_sum = local_pes_9_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_12_io_in_sum_exp = local_pes_9_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_12_io_in_kv = local_pes_8_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_12_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_12_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_12_io_in_stage = local_pes_9_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_13_clock = clock;
  assign local_pes_9_13_reset = reset;
  assign local_pes_9_13_io_in_q = local_pes_9_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_13_io_in_sum = local_pes_9_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_13_io_in_sum_exp = local_pes_9_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_13_io_in_kv = local_pes_8_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_13_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_13_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_13_io_in_stage = local_pes_9_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_14_clock = clock;
  assign local_pes_9_14_reset = reset;
  assign local_pes_9_14_io_in_q = local_pes_9_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_14_io_in_sum = local_pes_9_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_14_io_in_sum_exp = local_pes_9_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_14_io_in_kv = local_pes_8_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_14_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_14_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_14_io_in_stage = local_pes_9_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_15_clock = clock;
  assign local_pes_9_15_reset = reset;
  assign local_pes_9_15_io_in_q = local_pes_9_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_15_io_in_sum = local_pes_9_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_15_io_in_sum_exp = local_pes_9_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_15_io_in_kv = local_pes_8_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_15_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_15_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_15_io_in_stage = local_pes_9_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_16_clock = clock;
  assign local_pes_9_16_reset = reset;
  assign local_pes_9_16_io_in_q = local_pes_9_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_16_io_in_sum = local_pes_9_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_16_io_in_sum_exp = local_pes_9_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_16_io_in_kv = local_pes_8_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_16_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_16_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_16_io_in_stage = local_pes_9_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_17_clock = clock;
  assign local_pes_9_17_reset = reset;
  assign local_pes_9_17_io_in_q = local_pes_9_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_17_io_in_sum = local_pes_9_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_17_io_in_sum_exp = local_pes_9_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_17_io_in_kv = local_pes_8_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_17_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_17_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_17_io_in_stage = local_pes_9_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_18_clock = clock;
  assign local_pes_9_18_reset = reset;
  assign local_pes_9_18_io_in_q = local_pes_9_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_18_io_in_sum = local_pes_9_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_18_io_in_sum_exp = local_pes_9_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_18_io_in_kv = local_pes_8_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_18_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_18_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_18_io_in_stage = local_pes_9_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_19_clock = clock;
  assign local_pes_9_19_reset = reset;
  assign local_pes_9_19_io_in_q = local_pes_9_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_19_io_in_sum = local_pes_9_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_19_io_in_sum_exp = local_pes_9_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_19_io_in_kv = local_pes_8_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_19_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_19_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_19_io_in_stage = local_pes_9_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_20_clock = clock;
  assign local_pes_9_20_reset = reset;
  assign local_pes_9_20_io_in_q = local_pes_9_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_20_io_in_sum = local_pes_9_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_20_io_in_sum_exp = local_pes_9_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_20_io_in_kv = local_pes_8_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_20_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_20_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_20_io_in_stage = local_pes_9_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_21_clock = clock;
  assign local_pes_9_21_reset = reset;
  assign local_pes_9_21_io_in_q = local_pes_9_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_21_io_in_sum = local_pes_9_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_21_io_in_sum_exp = local_pes_9_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_21_io_in_kv = local_pes_8_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_21_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_21_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_21_io_in_stage = local_pes_9_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_22_clock = clock;
  assign local_pes_9_22_reset = reset;
  assign local_pes_9_22_io_in_q = local_pes_9_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_22_io_in_sum = local_pes_9_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_22_io_in_sum_exp = local_pes_9_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_22_io_in_kv = local_pes_8_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_22_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_22_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_22_io_in_stage = local_pes_9_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_23_clock = clock;
  assign local_pes_9_23_reset = reset;
  assign local_pes_9_23_io_in_q = local_pes_9_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_23_io_in_sum = local_pes_9_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_23_io_in_sum_exp = local_pes_9_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_23_io_in_kv = local_pes_8_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_23_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_23_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_23_io_in_stage = local_pes_9_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_24_clock = clock;
  assign local_pes_9_24_reset = reset;
  assign local_pes_9_24_io_in_q = local_pes_9_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_24_io_in_sum = local_pes_9_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_24_io_in_sum_exp = local_pes_9_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_24_io_in_kv = local_pes_8_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_24_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_24_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_24_io_in_stage = local_pes_9_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_25_clock = clock;
  assign local_pes_9_25_reset = reset;
  assign local_pes_9_25_io_in_q = local_pes_9_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_25_io_in_sum = local_pes_9_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_25_io_in_sum_exp = local_pes_9_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_25_io_in_kv = local_pes_8_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_25_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_25_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_25_io_in_stage = local_pes_9_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_26_clock = clock;
  assign local_pes_9_26_reset = reset;
  assign local_pes_9_26_io_in_q = local_pes_9_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_26_io_in_sum = local_pes_9_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_26_io_in_sum_exp = local_pes_9_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_26_io_in_kv = local_pes_8_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_26_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_26_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_26_io_in_stage = local_pes_9_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_27_clock = clock;
  assign local_pes_9_27_reset = reset;
  assign local_pes_9_27_io_in_q = local_pes_9_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_27_io_in_sum = local_pes_9_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_27_io_in_sum_exp = local_pes_9_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_27_io_in_kv = local_pes_8_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_27_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_27_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_27_io_in_stage = local_pes_9_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_28_clock = clock;
  assign local_pes_9_28_reset = reset;
  assign local_pes_9_28_io_in_q = local_pes_9_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_28_io_in_sum = local_pes_9_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_28_io_in_sum_exp = local_pes_9_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_28_io_in_kv = local_pes_8_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_28_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_28_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_28_io_in_stage = local_pes_9_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_29_clock = clock;
  assign local_pes_9_29_reset = reset;
  assign local_pes_9_29_io_in_q = local_pes_9_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_29_io_in_sum = local_pes_9_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_29_io_in_sum_exp = local_pes_9_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_29_io_in_kv = local_pes_8_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_29_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_29_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_29_io_in_stage = local_pes_9_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_30_clock = clock;
  assign local_pes_9_30_reset = reset;
  assign local_pes_9_30_io_in_q = local_pes_9_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_30_io_in_sum = local_pes_9_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_30_io_in_sum_exp = local_pes_9_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_30_io_in_kv = local_pes_8_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_30_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_30_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_30_io_in_stage = local_pes_9_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_9_31_clock = clock;
  assign local_pes_9_31_reset = reset;
  assign local_pes_9_31_io_in_q = local_pes_9_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_9_31_io_in_sum = local_pes_9_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_9_31_io_in_sum_exp = local_pes_9_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_9_31_io_in_kv = local_pes_8_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_9_31_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_9_31_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_9_31_io_in_stage = local_pes_9_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_0_clock = clock;
  assign local_pes_10_0_reset = reset;
  assign local_pes_10_0_io_in_q = io_q_ports_10; // @[PEArray.scala 51:37]
  assign local_pes_10_0_io_in_kv = io_kv_ports_41; // @[PEArray.scala 40:34]
  assign local_pes_10_0_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_0_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_0_io_in_stage = io_stage_ports_10; // @[PEArray.scala 52:41]
  assign local_pes_10_1_clock = clock;
  assign local_pes_10_1_reset = reset;
  assign local_pes_10_1_io_in_q = local_pes_10_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_1_io_in_sum = local_pes_10_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_10_1_io_in_kv = local_pes_9_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_1_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_1_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_1_io_in_stage = local_pes_10_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_2_clock = clock;
  assign local_pes_10_2_reset = reset;
  assign local_pes_10_2_io_in_q = local_pes_10_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_2_io_in_sum = local_pes_10_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_2_io_in_sum_exp = local_pes_10_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_2_io_in_kv = local_pes_9_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_2_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_2_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_2_io_in_stage = local_pes_10_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_3_clock = clock;
  assign local_pes_10_3_reset = reset;
  assign local_pes_10_3_io_in_q = local_pes_10_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_3_io_in_sum = local_pes_10_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_3_io_in_sum_exp = local_pes_10_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_3_io_in_kv = local_pes_9_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_3_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_3_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_3_io_in_stage = local_pes_10_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_4_clock = clock;
  assign local_pes_10_4_reset = reset;
  assign local_pes_10_4_io_in_q = local_pes_10_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_4_io_in_sum = local_pes_10_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_4_io_in_sum_exp = local_pes_10_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_4_io_in_kv = local_pes_9_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_4_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_4_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_4_io_in_stage = local_pes_10_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_5_clock = clock;
  assign local_pes_10_5_reset = reset;
  assign local_pes_10_5_io_in_q = local_pes_10_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_5_io_in_sum = local_pes_10_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_5_io_in_sum_exp = local_pes_10_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_5_io_in_kv = local_pes_9_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_5_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_5_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_5_io_in_stage = local_pes_10_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_6_clock = clock;
  assign local_pes_10_6_reset = reset;
  assign local_pes_10_6_io_in_q = local_pes_10_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_6_io_in_sum = local_pes_10_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_6_io_in_sum_exp = local_pes_10_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_6_io_in_kv = local_pes_9_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_6_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_6_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_6_io_in_stage = local_pes_10_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_7_clock = clock;
  assign local_pes_10_7_reset = reset;
  assign local_pes_10_7_io_in_q = local_pes_10_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_7_io_in_sum = local_pes_10_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_7_io_in_sum_exp = local_pes_10_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_7_io_in_kv = local_pes_9_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_7_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_7_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_7_io_in_stage = local_pes_10_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_8_clock = clock;
  assign local_pes_10_8_reset = reset;
  assign local_pes_10_8_io_in_q = local_pes_10_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_8_io_in_sum = local_pes_10_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_8_io_in_sum_exp = local_pes_10_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_8_io_in_kv = local_pes_9_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_8_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_8_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_8_io_in_stage = local_pes_10_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_9_clock = clock;
  assign local_pes_10_9_reset = reset;
  assign local_pes_10_9_io_in_q = local_pes_10_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_9_io_in_sum = local_pes_10_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_9_io_in_sum_exp = local_pes_10_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_9_io_in_kv = local_pes_9_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_9_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_9_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_9_io_in_stage = local_pes_10_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_10_clock = clock;
  assign local_pes_10_10_reset = reset;
  assign local_pes_10_10_io_in_q = local_pes_10_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_10_io_in_sum = local_pes_10_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_10_io_in_sum_exp = local_pes_10_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_10_io_in_kv = local_pes_9_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_10_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_10_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_10_io_in_stage = local_pes_10_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_11_clock = clock;
  assign local_pes_10_11_reset = reset;
  assign local_pes_10_11_io_in_q = local_pes_10_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_11_io_in_sum = local_pes_10_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_11_io_in_sum_exp = local_pes_10_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_11_io_in_kv = local_pes_9_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_11_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_11_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_11_io_in_stage = local_pes_10_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_12_clock = clock;
  assign local_pes_10_12_reset = reset;
  assign local_pes_10_12_io_in_q = local_pes_10_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_12_io_in_sum = local_pes_10_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_12_io_in_sum_exp = local_pes_10_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_12_io_in_kv = local_pes_9_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_12_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_12_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_12_io_in_stage = local_pes_10_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_13_clock = clock;
  assign local_pes_10_13_reset = reset;
  assign local_pes_10_13_io_in_q = local_pes_10_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_13_io_in_sum = local_pes_10_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_13_io_in_sum_exp = local_pes_10_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_13_io_in_kv = local_pes_9_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_13_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_13_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_13_io_in_stage = local_pes_10_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_14_clock = clock;
  assign local_pes_10_14_reset = reset;
  assign local_pes_10_14_io_in_q = local_pes_10_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_14_io_in_sum = local_pes_10_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_14_io_in_sum_exp = local_pes_10_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_14_io_in_kv = local_pes_9_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_14_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_14_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_14_io_in_stage = local_pes_10_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_15_clock = clock;
  assign local_pes_10_15_reset = reset;
  assign local_pes_10_15_io_in_q = local_pes_10_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_15_io_in_sum = local_pes_10_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_15_io_in_sum_exp = local_pes_10_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_15_io_in_kv = local_pes_9_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_15_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_15_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_15_io_in_stage = local_pes_10_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_16_clock = clock;
  assign local_pes_10_16_reset = reset;
  assign local_pes_10_16_io_in_q = local_pes_10_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_16_io_in_sum = local_pes_10_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_16_io_in_sum_exp = local_pes_10_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_16_io_in_kv = local_pes_9_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_16_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_16_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_16_io_in_stage = local_pes_10_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_17_clock = clock;
  assign local_pes_10_17_reset = reset;
  assign local_pes_10_17_io_in_q = local_pes_10_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_17_io_in_sum = local_pes_10_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_17_io_in_sum_exp = local_pes_10_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_17_io_in_kv = local_pes_9_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_17_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_17_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_17_io_in_stage = local_pes_10_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_18_clock = clock;
  assign local_pes_10_18_reset = reset;
  assign local_pes_10_18_io_in_q = local_pes_10_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_18_io_in_sum = local_pes_10_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_18_io_in_sum_exp = local_pes_10_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_18_io_in_kv = local_pes_9_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_18_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_18_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_18_io_in_stage = local_pes_10_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_19_clock = clock;
  assign local_pes_10_19_reset = reset;
  assign local_pes_10_19_io_in_q = local_pes_10_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_19_io_in_sum = local_pes_10_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_19_io_in_sum_exp = local_pes_10_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_19_io_in_kv = local_pes_9_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_19_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_19_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_19_io_in_stage = local_pes_10_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_20_clock = clock;
  assign local_pes_10_20_reset = reset;
  assign local_pes_10_20_io_in_q = local_pes_10_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_20_io_in_sum = local_pes_10_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_20_io_in_sum_exp = local_pes_10_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_20_io_in_kv = local_pes_9_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_20_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_20_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_20_io_in_stage = local_pes_10_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_21_clock = clock;
  assign local_pes_10_21_reset = reset;
  assign local_pes_10_21_io_in_q = local_pes_10_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_21_io_in_sum = local_pes_10_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_21_io_in_sum_exp = local_pes_10_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_21_io_in_kv = local_pes_9_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_21_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_21_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_21_io_in_stage = local_pes_10_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_22_clock = clock;
  assign local_pes_10_22_reset = reset;
  assign local_pes_10_22_io_in_q = local_pes_10_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_22_io_in_sum = local_pes_10_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_22_io_in_sum_exp = local_pes_10_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_22_io_in_kv = local_pes_9_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_22_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_22_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_22_io_in_stage = local_pes_10_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_23_clock = clock;
  assign local_pes_10_23_reset = reset;
  assign local_pes_10_23_io_in_q = local_pes_10_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_23_io_in_sum = local_pes_10_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_23_io_in_sum_exp = local_pes_10_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_23_io_in_kv = local_pes_9_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_23_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_23_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_23_io_in_stage = local_pes_10_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_24_clock = clock;
  assign local_pes_10_24_reset = reset;
  assign local_pes_10_24_io_in_q = local_pes_10_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_24_io_in_sum = local_pes_10_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_24_io_in_sum_exp = local_pes_10_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_24_io_in_kv = local_pes_9_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_24_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_24_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_24_io_in_stage = local_pes_10_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_25_clock = clock;
  assign local_pes_10_25_reset = reset;
  assign local_pes_10_25_io_in_q = local_pes_10_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_25_io_in_sum = local_pes_10_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_25_io_in_sum_exp = local_pes_10_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_25_io_in_kv = local_pes_9_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_25_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_25_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_25_io_in_stage = local_pes_10_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_26_clock = clock;
  assign local_pes_10_26_reset = reset;
  assign local_pes_10_26_io_in_q = local_pes_10_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_26_io_in_sum = local_pes_10_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_26_io_in_sum_exp = local_pes_10_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_26_io_in_kv = local_pes_9_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_26_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_26_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_26_io_in_stage = local_pes_10_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_27_clock = clock;
  assign local_pes_10_27_reset = reset;
  assign local_pes_10_27_io_in_q = local_pes_10_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_27_io_in_sum = local_pes_10_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_27_io_in_sum_exp = local_pes_10_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_27_io_in_kv = local_pes_9_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_27_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_27_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_27_io_in_stage = local_pes_10_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_28_clock = clock;
  assign local_pes_10_28_reset = reset;
  assign local_pes_10_28_io_in_q = local_pes_10_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_28_io_in_sum = local_pes_10_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_28_io_in_sum_exp = local_pes_10_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_28_io_in_kv = local_pes_9_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_28_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_28_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_28_io_in_stage = local_pes_10_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_29_clock = clock;
  assign local_pes_10_29_reset = reset;
  assign local_pes_10_29_io_in_q = local_pes_10_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_29_io_in_sum = local_pes_10_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_29_io_in_sum_exp = local_pes_10_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_29_io_in_kv = local_pes_9_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_29_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_29_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_29_io_in_stage = local_pes_10_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_30_clock = clock;
  assign local_pes_10_30_reset = reset;
  assign local_pes_10_30_io_in_q = local_pes_10_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_30_io_in_sum = local_pes_10_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_30_io_in_sum_exp = local_pes_10_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_30_io_in_kv = local_pes_9_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_30_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_30_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_30_io_in_stage = local_pes_10_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_10_31_clock = clock;
  assign local_pes_10_31_reset = reset;
  assign local_pes_10_31_io_in_q = local_pes_10_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_10_31_io_in_sum = local_pes_10_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_10_31_io_in_sum_exp = local_pes_10_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_10_31_io_in_kv = local_pes_9_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_10_31_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_10_31_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_10_31_io_in_stage = local_pes_10_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_0_clock = clock;
  assign local_pes_11_0_reset = reset;
  assign local_pes_11_0_io_in_q = io_q_ports_11; // @[PEArray.scala 51:37]
  assign local_pes_11_0_io_in_kv = io_kv_ports_42; // @[PEArray.scala 40:34]
  assign local_pes_11_0_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_0_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_0_io_in_stage = io_stage_ports_11; // @[PEArray.scala 52:41]
  assign local_pes_11_1_clock = clock;
  assign local_pes_11_1_reset = reset;
  assign local_pes_11_1_io_in_q = local_pes_11_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_1_io_in_sum = local_pes_11_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_11_1_io_in_kv = local_pes_10_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_1_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_1_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_1_io_in_stage = local_pes_11_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_2_clock = clock;
  assign local_pes_11_2_reset = reset;
  assign local_pes_11_2_io_in_q = local_pes_11_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_2_io_in_sum = local_pes_11_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_2_io_in_sum_exp = local_pes_11_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_2_io_in_kv = local_pes_10_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_2_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_2_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_2_io_in_stage = local_pes_11_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_3_clock = clock;
  assign local_pes_11_3_reset = reset;
  assign local_pes_11_3_io_in_q = local_pes_11_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_3_io_in_sum = local_pes_11_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_3_io_in_sum_exp = local_pes_11_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_3_io_in_kv = local_pes_10_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_3_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_3_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_3_io_in_stage = local_pes_11_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_4_clock = clock;
  assign local_pes_11_4_reset = reset;
  assign local_pes_11_4_io_in_q = local_pes_11_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_4_io_in_sum = local_pes_11_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_4_io_in_sum_exp = local_pes_11_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_4_io_in_kv = local_pes_10_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_4_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_4_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_4_io_in_stage = local_pes_11_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_5_clock = clock;
  assign local_pes_11_5_reset = reset;
  assign local_pes_11_5_io_in_q = local_pes_11_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_5_io_in_sum = local_pes_11_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_5_io_in_sum_exp = local_pes_11_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_5_io_in_kv = local_pes_10_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_5_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_5_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_5_io_in_stage = local_pes_11_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_6_clock = clock;
  assign local_pes_11_6_reset = reset;
  assign local_pes_11_6_io_in_q = local_pes_11_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_6_io_in_sum = local_pes_11_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_6_io_in_sum_exp = local_pes_11_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_6_io_in_kv = local_pes_10_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_6_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_6_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_6_io_in_stage = local_pes_11_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_7_clock = clock;
  assign local_pes_11_7_reset = reset;
  assign local_pes_11_7_io_in_q = local_pes_11_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_7_io_in_sum = local_pes_11_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_7_io_in_sum_exp = local_pes_11_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_7_io_in_kv = local_pes_10_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_7_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_7_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_7_io_in_stage = local_pes_11_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_8_clock = clock;
  assign local_pes_11_8_reset = reset;
  assign local_pes_11_8_io_in_q = local_pes_11_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_8_io_in_sum = local_pes_11_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_8_io_in_sum_exp = local_pes_11_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_8_io_in_kv = local_pes_10_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_8_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_8_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_8_io_in_stage = local_pes_11_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_9_clock = clock;
  assign local_pes_11_9_reset = reset;
  assign local_pes_11_9_io_in_q = local_pes_11_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_9_io_in_sum = local_pes_11_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_9_io_in_sum_exp = local_pes_11_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_9_io_in_kv = local_pes_10_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_9_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_9_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_9_io_in_stage = local_pes_11_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_10_clock = clock;
  assign local_pes_11_10_reset = reset;
  assign local_pes_11_10_io_in_q = local_pes_11_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_10_io_in_sum = local_pes_11_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_10_io_in_sum_exp = local_pes_11_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_10_io_in_kv = local_pes_10_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_10_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_10_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_10_io_in_stage = local_pes_11_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_11_clock = clock;
  assign local_pes_11_11_reset = reset;
  assign local_pes_11_11_io_in_q = local_pes_11_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_11_io_in_sum = local_pes_11_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_11_io_in_sum_exp = local_pes_11_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_11_io_in_kv = local_pes_10_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_11_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_11_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_11_io_in_stage = local_pes_11_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_12_clock = clock;
  assign local_pes_11_12_reset = reset;
  assign local_pes_11_12_io_in_q = local_pes_11_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_12_io_in_sum = local_pes_11_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_12_io_in_sum_exp = local_pes_11_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_12_io_in_kv = local_pes_10_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_12_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_12_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_12_io_in_stage = local_pes_11_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_13_clock = clock;
  assign local_pes_11_13_reset = reset;
  assign local_pes_11_13_io_in_q = local_pes_11_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_13_io_in_sum = local_pes_11_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_13_io_in_sum_exp = local_pes_11_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_13_io_in_kv = local_pes_10_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_13_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_13_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_13_io_in_stage = local_pes_11_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_14_clock = clock;
  assign local_pes_11_14_reset = reset;
  assign local_pes_11_14_io_in_q = local_pes_11_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_14_io_in_sum = local_pes_11_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_14_io_in_sum_exp = local_pes_11_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_14_io_in_kv = local_pes_10_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_14_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_14_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_14_io_in_stage = local_pes_11_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_15_clock = clock;
  assign local_pes_11_15_reset = reset;
  assign local_pes_11_15_io_in_q = local_pes_11_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_15_io_in_sum = local_pes_11_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_15_io_in_sum_exp = local_pes_11_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_15_io_in_kv = local_pes_10_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_15_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_15_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_15_io_in_stage = local_pes_11_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_16_clock = clock;
  assign local_pes_11_16_reset = reset;
  assign local_pes_11_16_io_in_q = local_pes_11_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_16_io_in_sum = local_pes_11_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_16_io_in_sum_exp = local_pes_11_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_16_io_in_kv = local_pes_10_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_16_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_16_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_16_io_in_stage = local_pes_11_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_17_clock = clock;
  assign local_pes_11_17_reset = reset;
  assign local_pes_11_17_io_in_q = local_pes_11_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_17_io_in_sum = local_pes_11_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_17_io_in_sum_exp = local_pes_11_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_17_io_in_kv = local_pes_10_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_17_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_17_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_17_io_in_stage = local_pes_11_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_18_clock = clock;
  assign local_pes_11_18_reset = reset;
  assign local_pes_11_18_io_in_q = local_pes_11_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_18_io_in_sum = local_pes_11_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_18_io_in_sum_exp = local_pes_11_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_18_io_in_kv = local_pes_10_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_18_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_18_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_18_io_in_stage = local_pes_11_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_19_clock = clock;
  assign local_pes_11_19_reset = reset;
  assign local_pes_11_19_io_in_q = local_pes_11_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_19_io_in_sum = local_pes_11_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_19_io_in_sum_exp = local_pes_11_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_19_io_in_kv = local_pes_10_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_19_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_19_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_19_io_in_stage = local_pes_11_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_20_clock = clock;
  assign local_pes_11_20_reset = reset;
  assign local_pes_11_20_io_in_q = local_pes_11_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_20_io_in_sum = local_pes_11_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_20_io_in_sum_exp = local_pes_11_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_20_io_in_kv = local_pes_10_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_20_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_20_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_20_io_in_stage = local_pes_11_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_21_clock = clock;
  assign local_pes_11_21_reset = reset;
  assign local_pes_11_21_io_in_q = local_pes_11_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_21_io_in_sum = local_pes_11_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_21_io_in_sum_exp = local_pes_11_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_21_io_in_kv = local_pes_10_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_21_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_21_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_21_io_in_stage = local_pes_11_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_22_clock = clock;
  assign local_pes_11_22_reset = reset;
  assign local_pes_11_22_io_in_q = local_pes_11_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_22_io_in_sum = local_pes_11_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_22_io_in_sum_exp = local_pes_11_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_22_io_in_kv = local_pes_10_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_22_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_22_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_22_io_in_stage = local_pes_11_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_23_clock = clock;
  assign local_pes_11_23_reset = reset;
  assign local_pes_11_23_io_in_q = local_pes_11_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_23_io_in_sum = local_pes_11_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_23_io_in_sum_exp = local_pes_11_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_23_io_in_kv = local_pes_10_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_23_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_23_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_23_io_in_stage = local_pes_11_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_24_clock = clock;
  assign local_pes_11_24_reset = reset;
  assign local_pes_11_24_io_in_q = local_pes_11_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_24_io_in_sum = local_pes_11_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_24_io_in_sum_exp = local_pes_11_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_24_io_in_kv = local_pes_10_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_24_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_24_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_24_io_in_stage = local_pes_11_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_25_clock = clock;
  assign local_pes_11_25_reset = reset;
  assign local_pes_11_25_io_in_q = local_pes_11_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_25_io_in_sum = local_pes_11_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_25_io_in_sum_exp = local_pes_11_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_25_io_in_kv = local_pes_10_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_25_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_25_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_25_io_in_stage = local_pes_11_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_26_clock = clock;
  assign local_pes_11_26_reset = reset;
  assign local_pes_11_26_io_in_q = local_pes_11_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_26_io_in_sum = local_pes_11_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_26_io_in_sum_exp = local_pes_11_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_26_io_in_kv = local_pes_10_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_26_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_26_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_26_io_in_stage = local_pes_11_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_27_clock = clock;
  assign local_pes_11_27_reset = reset;
  assign local_pes_11_27_io_in_q = local_pes_11_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_27_io_in_sum = local_pes_11_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_27_io_in_sum_exp = local_pes_11_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_27_io_in_kv = local_pes_10_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_27_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_27_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_27_io_in_stage = local_pes_11_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_28_clock = clock;
  assign local_pes_11_28_reset = reset;
  assign local_pes_11_28_io_in_q = local_pes_11_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_28_io_in_sum = local_pes_11_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_28_io_in_sum_exp = local_pes_11_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_28_io_in_kv = local_pes_10_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_28_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_28_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_28_io_in_stage = local_pes_11_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_29_clock = clock;
  assign local_pes_11_29_reset = reset;
  assign local_pes_11_29_io_in_q = local_pes_11_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_29_io_in_sum = local_pes_11_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_29_io_in_sum_exp = local_pes_11_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_29_io_in_kv = local_pes_10_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_29_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_29_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_29_io_in_stage = local_pes_11_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_30_clock = clock;
  assign local_pes_11_30_reset = reset;
  assign local_pes_11_30_io_in_q = local_pes_11_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_30_io_in_sum = local_pes_11_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_30_io_in_sum_exp = local_pes_11_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_30_io_in_kv = local_pes_10_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_30_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_30_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_30_io_in_stage = local_pes_11_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_11_31_clock = clock;
  assign local_pes_11_31_reset = reset;
  assign local_pes_11_31_io_in_q = local_pes_11_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_11_31_io_in_sum = local_pes_11_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_11_31_io_in_sum_exp = local_pes_11_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_11_31_io_in_kv = local_pes_10_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_11_31_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_11_31_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_11_31_io_in_stage = local_pes_11_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_0_clock = clock;
  assign local_pes_12_0_reset = reset;
  assign local_pes_12_0_io_in_q = io_q_ports_12; // @[PEArray.scala 51:37]
  assign local_pes_12_0_io_in_kv = io_kv_ports_43; // @[PEArray.scala 40:34]
  assign local_pes_12_0_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_0_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_0_io_in_stage = io_stage_ports_12; // @[PEArray.scala 52:41]
  assign local_pes_12_1_clock = clock;
  assign local_pes_12_1_reset = reset;
  assign local_pes_12_1_io_in_q = local_pes_12_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_1_io_in_sum = local_pes_12_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_12_1_io_in_kv = local_pes_11_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_1_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_1_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_1_io_in_stage = local_pes_12_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_2_clock = clock;
  assign local_pes_12_2_reset = reset;
  assign local_pes_12_2_io_in_q = local_pes_12_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_2_io_in_sum = local_pes_12_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_2_io_in_sum_exp = local_pes_12_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_2_io_in_kv = local_pes_11_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_2_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_2_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_2_io_in_stage = local_pes_12_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_3_clock = clock;
  assign local_pes_12_3_reset = reset;
  assign local_pes_12_3_io_in_q = local_pes_12_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_3_io_in_sum = local_pes_12_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_3_io_in_sum_exp = local_pes_12_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_3_io_in_kv = local_pes_11_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_3_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_3_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_3_io_in_stage = local_pes_12_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_4_clock = clock;
  assign local_pes_12_4_reset = reset;
  assign local_pes_12_4_io_in_q = local_pes_12_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_4_io_in_sum = local_pes_12_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_4_io_in_sum_exp = local_pes_12_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_4_io_in_kv = local_pes_11_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_4_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_4_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_4_io_in_stage = local_pes_12_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_5_clock = clock;
  assign local_pes_12_5_reset = reset;
  assign local_pes_12_5_io_in_q = local_pes_12_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_5_io_in_sum = local_pes_12_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_5_io_in_sum_exp = local_pes_12_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_5_io_in_kv = local_pes_11_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_5_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_5_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_5_io_in_stage = local_pes_12_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_6_clock = clock;
  assign local_pes_12_6_reset = reset;
  assign local_pes_12_6_io_in_q = local_pes_12_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_6_io_in_sum = local_pes_12_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_6_io_in_sum_exp = local_pes_12_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_6_io_in_kv = local_pes_11_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_6_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_6_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_6_io_in_stage = local_pes_12_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_7_clock = clock;
  assign local_pes_12_7_reset = reset;
  assign local_pes_12_7_io_in_q = local_pes_12_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_7_io_in_sum = local_pes_12_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_7_io_in_sum_exp = local_pes_12_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_7_io_in_kv = local_pes_11_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_7_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_7_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_7_io_in_stage = local_pes_12_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_8_clock = clock;
  assign local_pes_12_8_reset = reset;
  assign local_pes_12_8_io_in_q = local_pes_12_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_8_io_in_sum = local_pes_12_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_8_io_in_sum_exp = local_pes_12_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_8_io_in_kv = local_pes_11_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_8_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_8_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_8_io_in_stage = local_pes_12_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_9_clock = clock;
  assign local_pes_12_9_reset = reset;
  assign local_pes_12_9_io_in_q = local_pes_12_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_9_io_in_sum = local_pes_12_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_9_io_in_sum_exp = local_pes_12_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_9_io_in_kv = local_pes_11_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_9_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_9_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_9_io_in_stage = local_pes_12_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_10_clock = clock;
  assign local_pes_12_10_reset = reset;
  assign local_pes_12_10_io_in_q = local_pes_12_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_10_io_in_sum = local_pes_12_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_10_io_in_sum_exp = local_pes_12_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_10_io_in_kv = local_pes_11_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_10_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_10_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_10_io_in_stage = local_pes_12_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_11_clock = clock;
  assign local_pes_12_11_reset = reset;
  assign local_pes_12_11_io_in_q = local_pes_12_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_11_io_in_sum = local_pes_12_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_11_io_in_sum_exp = local_pes_12_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_11_io_in_kv = local_pes_11_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_11_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_11_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_11_io_in_stage = local_pes_12_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_12_clock = clock;
  assign local_pes_12_12_reset = reset;
  assign local_pes_12_12_io_in_q = local_pes_12_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_12_io_in_sum = local_pes_12_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_12_io_in_sum_exp = local_pes_12_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_12_io_in_kv = local_pes_11_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_12_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_12_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_12_io_in_stage = local_pes_12_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_13_clock = clock;
  assign local_pes_12_13_reset = reset;
  assign local_pes_12_13_io_in_q = local_pes_12_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_13_io_in_sum = local_pes_12_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_13_io_in_sum_exp = local_pes_12_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_13_io_in_kv = local_pes_11_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_13_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_13_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_13_io_in_stage = local_pes_12_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_14_clock = clock;
  assign local_pes_12_14_reset = reset;
  assign local_pes_12_14_io_in_q = local_pes_12_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_14_io_in_sum = local_pes_12_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_14_io_in_sum_exp = local_pes_12_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_14_io_in_kv = local_pes_11_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_14_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_14_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_14_io_in_stage = local_pes_12_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_15_clock = clock;
  assign local_pes_12_15_reset = reset;
  assign local_pes_12_15_io_in_q = local_pes_12_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_15_io_in_sum = local_pes_12_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_15_io_in_sum_exp = local_pes_12_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_15_io_in_kv = local_pes_11_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_15_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_15_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_15_io_in_stage = local_pes_12_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_16_clock = clock;
  assign local_pes_12_16_reset = reset;
  assign local_pes_12_16_io_in_q = local_pes_12_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_16_io_in_sum = local_pes_12_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_16_io_in_sum_exp = local_pes_12_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_16_io_in_kv = local_pes_11_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_16_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_16_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_16_io_in_stage = local_pes_12_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_17_clock = clock;
  assign local_pes_12_17_reset = reset;
  assign local_pes_12_17_io_in_q = local_pes_12_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_17_io_in_sum = local_pes_12_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_17_io_in_sum_exp = local_pes_12_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_17_io_in_kv = local_pes_11_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_17_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_17_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_17_io_in_stage = local_pes_12_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_18_clock = clock;
  assign local_pes_12_18_reset = reset;
  assign local_pes_12_18_io_in_q = local_pes_12_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_18_io_in_sum = local_pes_12_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_18_io_in_sum_exp = local_pes_12_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_18_io_in_kv = local_pes_11_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_18_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_18_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_18_io_in_stage = local_pes_12_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_19_clock = clock;
  assign local_pes_12_19_reset = reset;
  assign local_pes_12_19_io_in_q = local_pes_12_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_19_io_in_sum = local_pes_12_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_19_io_in_sum_exp = local_pes_12_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_19_io_in_kv = local_pes_11_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_19_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_19_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_19_io_in_stage = local_pes_12_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_20_clock = clock;
  assign local_pes_12_20_reset = reset;
  assign local_pes_12_20_io_in_q = local_pes_12_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_20_io_in_sum = local_pes_12_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_20_io_in_sum_exp = local_pes_12_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_20_io_in_kv = local_pes_11_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_20_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_20_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_20_io_in_stage = local_pes_12_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_21_clock = clock;
  assign local_pes_12_21_reset = reset;
  assign local_pes_12_21_io_in_q = local_pes_12_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_21_io_in_sum = local_pes_12_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_21_io_in_sum_exp = local_pes_12_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_21_io_in_kv = local_pes_11_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_21_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_21_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_21_io_in_stage = local_pes_12_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_22_clock = clock;
  assign local_pes_12_22_reset = reset;
  assign local_pes_12_22_io_in_q = local_pes_12_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_22_io_in_sum = local_pes_12_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_22_io_in_sum_exp = local_pes_12_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_22_io_in_kv = local_pes_11_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_22_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_22_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_22_io_in_stage = local_pes_12_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_23_clock = clock;
  assign local_pes_12_23_reset = reset;
  assign local_pes_12_23_io_in_q = local_pes_12_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_23_io_in_sum = local_pes_12_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_23_io_in_sum_exp = local_pes_12_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_23_io_in_kv = local_pes_11_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_23_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_23_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_23_io_in_stage = local_pes_12_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_24_clock = clock;
  assign local_pes_12_24_reset = reset;
  assign local_pes_12_24_io_in_q = local_pes_12_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_24_io_in_sum = local_pes_12_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_24_io_in_sum_exp = local_pes_12_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_24_io_in_kv = local_pes_11_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_24_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_24_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_24_io_in_stage = local_pes_12_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_25_clock = clock;
  assign local_pes_12_25_reset = reset;
  assign local_pes_12_25_io_in_q = local_pes_12_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_25_io_in_sum = local_pes_12_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_25_io_in_sum_exp = local_pes_12_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_25_io_in_kv = local_pes_11_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_25_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_25_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_25_io_in_stage = local_pes_12_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_26_clock = clock;
  assign local_pes_12_26_reset = reset;
  assign local_pes_12_26_io_in_q = local_pes_12_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_26_io_in_sum = local_pes_12_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_26_io_in_sum_exp = local_pes_12_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_26_io_in_kv = local_pes_11_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_26_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_26_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_26_io_in_stage = local_pes_12_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_27_clock = clock;
  assign local_pes_12_27_reset = reset;
  assign local_pes_12_27_io_in_q = local_pes_12_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_27_io_in_sum = local_pes_12_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_27_io_in_sum_exp = local_pes_12_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_27_io_in_kv = local_pes_11_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_27_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_27_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_27_io_in_stage = local_pes_12_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_28_clock = clock;
  assign local_pes_12_28_reset = reset;
  assign local_pes_12_28_io_in_q = local_pes_12_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_28_io_in_sum = local_pes_12_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_28_io_in_sum_exp = local_pes_12_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_28_io_in_kv = local_pes_11_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_28_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_28_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_28_io_in_stage = local_pes_12_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_29_clock = clock;
  assign local_pes_12_29_reset = reset;
  assign local_pes_12_29_io_in_q = local_pes_12_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_29_io_in_sum = local_pes_12_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_29_io_in_sum_exp = local_pes_12_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_29_io_in_kv = local_pes_11_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_29_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_29_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_29_io_in_stage = local_pes_12_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_30_clock = clock;
  assign local_pes_12_30_reset = reset;
  assign local_pes_12_30_io_in_q = local_pes_12_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_30_io_in_sum = local_pes_12_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_30_io_in_sum_exp = local_pes_12_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_30_io_in_kv = local_pes_11_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_30_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_30_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_30_io_in_stage = local_pes_12_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_12_31_clock = clock;
  assign local_pes_12_31_reset = reset;
  assign local_pes_12_31_io_in_q = local_pes_12_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_12_31_io_in_sum = local_pes_12_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_12_31_io_in_sum_exp = local_pes_12_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_12_31_io_in_kv = local_pes_11_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_12_31_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_12_31_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_12_31_io_in_stage = local_pes_12_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_0_clock = clock;
  assign local_pes_13_0_reset = reset;
  assign local_pes_13_0_io_in_q = io_q_ports_13; // @[PEArray.scala 51:37]
  assign local_pes_13_0_io_in_kv = io_kv_ports_44; // @[PEArray.scala 40:34]
  assign local_pes_13_0_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_0_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_0_io_in_stage = io_stage_ports_13; // @[PEArray.scala 52:41]
  assign local_pes_13_1_clock = clock;
  assign local_pes_13_1_reset = reset;
  assign local_pes_13_1_io_in_q = local_pes_13_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_1_io_in_sum = local_pes_13_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_13_1_io_in_kv = local_pes_12_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_1_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_1_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_1_io_in_stage = local_pes_13_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_2_clock = clock;
  assign local_pes_13_2_reset = reset;
  assign local_pes_13_2_io_in_q = local_pes_13_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_2_io_in_sum = local_pes_13_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_2_io_in_sum_exp = local_pes_13_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_2_io_in_kv = local_pes_12_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_2_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_2_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_2_io_in_stage = local_pes_13_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_3_clock = clock;
  assign local_pes_13_3_reset = reset;
  assign local_pes_13_3_io_in_q = local_pes_13_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_3_io_in_sum = local_pes_13_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_3_io_in_sum_exp = local_pes_13_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_3_io_in_kv = local_pes_12_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_3_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_3_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_3_io_in_stage = local_pes_13_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_4_clock = clock;
  assign local_pes_13_4_reset = reset;
  assign local_pes_13_4_io_in_q = local_pes_13_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_4_io_in_sum = local_pes_13_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_4_io_in_sum_exp = local_pes_13_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_4_io_in_kv = local_pes_12_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_4_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_4_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_4_io_in_stage = local_pes_13_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_5_clock = clock;
  assign local_pes_13_5_reset = reset;
  assign local_pes_13_5_io_in_q = local_pes_13_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_5_io_in_sum = local_pes_13_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_5_io_in_sum_exp = local_pes_13_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_5_io_in_kv = local_pes_12_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_5_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_5_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_5_io_in_stage = local_pes_13_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_6_clock = clock;
  assign local_pes_13_6_reset = reset;
  assign local_pes_13_6_io_in_q = local_pes_13_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_6_io_in_sum = local_pes_13_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_6_io_in_sum_exp = local_pes_13_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_6_io_in_kv = local_pes_12_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_6_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_6_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_6_io_in_stage = local_pes_13_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_7_clock = clock;
  assign local_pes_13_7_reset = reset;
  assign local_pes_13_7_io_in_q = local_pes_13_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_7_io_in_sum = local_pes_13_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_7_io_in_sum_exp = local_pes_13_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_7_io_in_kv = local_pes_12_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_7_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_7_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_7_io_in_stage = local_pes_13_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_8_clock = clock;
  assign local_pes_13_8_reset = reset;
  assign local_pes_13_8_io_in_q = local_pes_13_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_8_io_in_sum = local_pes_13_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_8_io_in_sum_exp = local_pes_13_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_8_io_in_kv = local_pes_12_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_8_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_8_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_8_io_in_stage = local_pes_13_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_9_clock = clock;
  assign local_pes_13_9_reset = reset;
  assign local_pes_13_9_io_in_q = local_pes_13_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_9_io_in_sum = local_pes_13_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_9_io_in_sum_exp = local_pes_13_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_9_io_in_kv = local_pes_12_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_9_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_9_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_9_io_in_stage = local_pes_13_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_10_clock = clock;
  assign local_pes_13_10_reset = reset;
  assign local_pes_13_10_io_in_q = local_pes_13_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_10_io_in_sum = local_pes_13_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_10_io_in_sum_exp = local_pes_13_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_10_io_in_kv = local_pes_12_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_10_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_10_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_10_io_in_stage = local_pes_13_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_11_clock = clock;
  assign local_pes_13_11_reset = reset;
  assign local_pes_13_11_io_in_q = local_pes_13_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_11_io_in_sum = local_pes_13_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_11_io_in_sum_exp = local_pes_13_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_11_io_in_kv = local_pes_12_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_11_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_11_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_11_io_in_stage = local_pes_13_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_12_clock = clock;
  assign local_pes_13_12_reset = reset;
  assign local_pes_13_12_io_in_q = local_pes_13_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_12_io_in_sum = local_pes_13_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_12_io_in_sum_exp = local_pes_13_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_12_io_in_kv = local_pes_12_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_12_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_12_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_12_io_in_stage = local_pes_13_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_13_clock = clock;
  assign local_pes_13_13_reset = reset;
  assign local_pes_13_13_io_in_q = local_pes_13_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_13_io_in_sum = local_pes_13_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_13_io_in_sum_exp = local_pes_13_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_13_io_in_kv = local_pes_12_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_13_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_13_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_13_io_in_stage = local_pes_13_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_14_clock = clock;
  assign local_pes_13_14_reset = reset;
  assign local_pes_13_14_io_in_q = local_pes_13_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_14_io_in_sum = local_pes_13_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_14_io_in_sum_exp = local_pes_13_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_14_io_in_kv = local_pes_12_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_14_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_14_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_14_io_in_stage = local_pes_13_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_15_clock = clock;
  assign local_pes_13_15_reset = reset;
  assign local_pes_13_15_io_in_q = local_pes_13_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_15_io_in_sum = local_pes_13_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_15_io_in_sum_exp = local_pes_13_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_15_io_in_kv = local_pes_12_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_15_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_15_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_15_io_in_stage = local_pes_13_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_16_clock = clock;
  assign local_pes_13_16_reset = reset;
  assign local_pes_13_16_io_in_q = local_pes_13_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_16_io_in_sum = local_pes_13_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_16_io_in_sum_exp = local_pes_13_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_16_io_in_kv = local_pes_12_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_16_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_16_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_16_io_in_stage = local_pes_13_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_17_clock = clock;
  assign local_pes_13_17_reset = reset;
  assign local_pes_13_17_io_in_q = local_pes_13_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_17_io_in_sum = local_pes_13_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_17_io_in_sum_exp = local_pes_13_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_17_io_in_kv = local_pes_12_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_17_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_17_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_17_io_in_stage = local_pes_13_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_18_clock = clock;
  assign local_pes_13_18_reset = reset;
  assign local_pes_13_18_io_in_q = local_pes_13_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_18_io_in_sum = local_pes_13_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_18_io_in_sum_exp = local_pes_13_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_18_io_in_kv = local_pes_12_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_18_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_18_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_18_io_in_stage = local_pes_13_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_19_clock = clock;
  assign local_pes_13_19_reset = reset;
  assign local_pes_13_19_io_in_q = local_pes_13_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_19_io_in_sum = local_pes_13_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_19_io_in_sum_exp = local_pes_13_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_19_io_in_kv = local_pes_12_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_19_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_19_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_19_io_in_stage = local_pes_13_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_20_clock = clock;
  assign local_pes_13_20_reset = reset;
  assign local_pes_13_20_io_in_q = local_pes_13_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_20_io_in_sum = local_pes_13_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_20_io_in_sum_exp = local_pes_13_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_20_io_in_kv = local_pes_12_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_20_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_20_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_20_io_in_stage = local_pes_13_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_21_clock = clock;
  assign local_pes_13_21_reset = reset;
  assign local_pes_13_21_io_in_q = local_pes_13_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_21_io_in_sum = local_pes_13_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_21_io_in_sum_exp = local_pes_13_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_21_io_in_kv = local_pes_12_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_21_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_21_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_21_io_in_stage = local_pes_13_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_22_clock = clock;
  assign local_pes_13_22_reset = reset;
  assign local_pes_13_22_io_in_q = local_pes_13_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_22_io_in_sum = local_pes_13_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_22_io_in_sum_exp = local_pes_13_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_22_io_in_kv = local_pes_12_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_22_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_22_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_22_io_in_stage = local_pes_13_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_23_clock = clock;
  assign local_pes_13_23_reset = reset;
  assign local_pes_13_23_io_in_q = local_pes_13_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_23_io_in_sum = local_pes_13_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_23_io_in_sum_exp = local_pes_13_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_23_io_in_kv = local_pes_12_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_23_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_23_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_23_io_in_stage = local_pes_13_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_24_clock = clock;
  assign local_pes_13_24_reset = reset;
  assign local_pes_13_24_io_in_q = local_pes_13_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_24_io_in_sum = local_pes_13_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_24_io_in_sum_exp = local_pes_13_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_24_io_in_kv = local_pes_12_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_24_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_24_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_24_io_in_stage = local_pes_13_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_25_clock = clock;
  assign local_pes_13_25_reset = reset;
  assign local_pes_13_25_io_in_q = local_pes_13_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_25_io_in_sum = local_pes_13_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_25_io_in_sum_exp = local_pes_13_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_25_io_in_kv = local_pes_12_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_25_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_25_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_25_io_in_stage = local_pes_13_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_26_clock = clock;
  assign local_pes_13_26_reset = reset;
  assign local_pes_13_26_io_in_q = local_pes_13_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_26_io_in_sum = local_pes_13_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_26_io_in_sum_exp = local_pes_13_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_26_io_in_kv = local_pes_12_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_26_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_26_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_26_io_in_stage = local_pes_13_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_27_clock = clock;
  assign local_pes_13_27_reset = reset;
  assign local_pes_13_27_io_in_q = local_pes_13_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_27_io_in_sum = local_pes_13_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_27_io_in_sum_exp = local_pes_13_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_27_io_in_kv = local_pes_12_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_27_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_27_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_27_io_in_stage = local_pes_13_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_28_clock = clock;
  assign local_pes_13_28_reset = reset;
  assign local_pes_13_28_io_in_q = local_pes_13_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_28_io_in_sum = local_pes_13_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_28_io_in_sum_exp = local_pes_13_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_28_io_in_kv = local_pes_12_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_28_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_28_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_28_io_in_stage = local_pes_13_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_29_clock = clock;
  assign local_pes_13_29_reset = reset;
  assign local_pes_13_29_io_in_q = local_pes_13_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_29_io_in_sum = local_pes_13_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_29_io_in_sum_exp = local_pes_13_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_29_io_in_kv = local_pes_12_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_29_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_29_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_29_io_in_stage = local_pes_13_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_30_clock = clock;
  assign local_pes_13_30_reset = reset;
  assign local_pes_13_30_io_in_q = local_pes_13_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_30_io_in_sum = local_pes_13_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_30_io_in_sum_exp = local_pes_13_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_30_io_in_kv = local_pes_12_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_30_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_30_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_30_io_in_stage = local_pes_13_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_13_31_clock = clock;
  assign local_pes_13_31_reset = reset;
  assign local_pes_13_31_io_in_q = local_pes_13_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_13_31_io_in_sum = local_pes_13_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_13_31_io_in_sum_exp = local_pes_13_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_13_31_io_in_kv = local_pes_12_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_13_31_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_13_31_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_13_31_io_in_stage = local_pes_13_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_0_clock = clock;
  assign local_pes_14_0_reset = reset;
  assign local_pes_14_0_io_in_q = io_q_ports_14; // @[PEArray.scala 51:37]
  assign local_pes_14_0_io_in_kv = io_kv_ports_45; // @[PEArray.scala 40:34]
  assign local_pes_14_0_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_0_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_0_io_in_stage = io_stage_ports_14; // @[PEArray.scala 52:41]
  assign local_pes_14_1_clock = clock;
  assign local_pes_14_1_reset = reset;
  assign local_pes_14_1_io_in_q = local_pes_14_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_1_io_in_sum = local_pes_14_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_14_1_io_in_kv = local_pes_13_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_1_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_1_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_1_io_in_stage = local_pes_14_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_2_clock = clock;
  assign local_pes_14_2_reset = reset;
  assign local_pes_14_2_io_in_q = local_pes_14_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_2_io_in_sum = local_pes_14_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_2_io_in_sum_exp = local_pes_14_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_2_io_in_kv = local_pes_13_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_2_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_2_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_2_io_in_stage = local_pes_14_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_3_clock = clock;
  assign local_pes_14_3_reset = reset;
  assign local_pes_14_3_io_in_q = local_pes_14_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_3_io_in_sum = local_pes_14_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_3_io_in_sum_exp = local_pes_14_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_3_io_in_kv = local_pes_13_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_3_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_3_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_3_io_in_stage = local_pes_14_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_4_clock = clock;
  assign local_pes_14_4_reset = reset;
  assign local_pes_14_4_io_in_q = local_pes_14_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_4_io_in_sum = local_pes_14_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_4_io_in_sum_exp = local_pes_14_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_4_io_in_kv = local_pes_13_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_4_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_4_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_4_io_in_stage = local_pes_14_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_5_clock = clock;
  assign local_pes_14_5_reset = reset;
  assign local_pes_14_5_io_in_q = local_pes_14_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_5_io_in_sum = local_pes_14_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_5_io_in_sum_exp = local_pes_14_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_5_io_in_kv = local_pes_13_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_5_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_5_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_5_io_in_stage = local_pes_14_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_6_clock = clock;
  assign local_pes_14_6_reset = reset;
  assign local_pes_14_6_io_in_q = local_pes_14_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_6_io_in_sum = local_pes_14_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_6_io_in_sum_exp = local_pes_14_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_6_io_in_kv = local_pes_13_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_6_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_6_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_6_io_in_stage = local_pes_14_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_7_clock = clock;
  assign local_pes_14_7_reset = reset;
  assign local_pes_14_7_io_in_q = local_pes_14_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_7_io_in_sum = local_pes_14_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_7_io_in_sum_exp = local_pes_14_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_7_io_in_kv = local_pes_13_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_7_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_7_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_7_io_in_stage = local_pes_14_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_8_clock = clock;
  assign local_pes_14_8_reset = reset;
  assign local_pes_14_8_io_in_q = local_pes_14_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_8_io_in_sum = local_pes_14_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_8_io_in_sum_exp = local_pes_14_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_8_io_in_kv = local_pes_13_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_8_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_8_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_8_io_in_stage = local_pes_14_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_9_clock = clock;
  assign local_pes_14_9_reset = reset;
  assign local_pes_14_9_io_in_q = local_pes_14_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_9_io_in_sum = local_pes_14_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_9_io_in_sum_exp = local_pes_14_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_9_io_in_kv = local_pes_13_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_9_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_9_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_9_io_in_stage = local_pes_14_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_10_clock = clock;
  assign local_pes_14_10_reset = reset;
  assign local_pes_14_10_io_in_q = local_pes_14_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_10_io_in_sum = local_pes_14_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_10_io_in_sum_exp = local_pes_14_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_10_io_in_kv = local_pes_13_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_10_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_10_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_10_io_in_stage = local_pes_14_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_11_clock = clock;
  assign local_pes_14_11_reset = reset;
  assign local_pes_14_11_io_in_q = local_pes_14_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_11_io_in_sum = local_pes_14_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_11_io_in_sum_exp = local_pes_14_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_11_io_in_kv = local_pes_13_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_11_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_11_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_11_io_in_stage = local_pes_14_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_12_clock = clock;
  assign local_pes_14_12_reset = reset;
  assign local_pes_14_12_io_in_q = local_pes_14_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_12_io_in_sum = local_pes_14_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_12_io_in_sum_exp = local_pes_14_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_12_io_in_kv = local_pes_13_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_12_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_12_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_12_io_in_stage = local_pes_14_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_13_clock = clock;
  assign local_pes_14_13_reset = reset;
  assign local_pes_14_13_io_in_q = local_pes_14_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_13_io_in_sum = local_pes_14_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_13_io_in_sum_exp = local_pes_14_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_13_io_in_kv = local_pes_13_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_13_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_13_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_13_io_in_stage = local_pes_14_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_14_clock = clock;
  assign local_pes_14_14_reset = reset;
  assign local_pes_14_14_io_in_q = local_pes_14_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_14_io_in_sum = local_pes_14_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_14_io_in_sum_exp = local_pes_14_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_14_io_in_kv = local_pes_13_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_14_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_14_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_14_io_in_stage = local_pes_14_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_15_clock = clock;
  assign local_pes_14_15_reset = reset;
  assign local_pes_14_15_io_in_q = local_pes_14_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_15_io_in_sum = local_pes_14_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_15_io_in_sum_exp = local_pes_14_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_15_io_in_kv = local_pes_13_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_15_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_15_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_15_io_in_stage = local_pes_14_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_16_clock = clock;
  assign local_pes_14_16_reset = reset;
  assign local_pes_14_16_io_in_q = local_pes_14_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_16_io_in_sum = local_pes_14_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_16_io_in_sum_exp = local_pes_14_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_16_io_in_kv = local_pes_13_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_16_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_16_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_16_io_in_stage = local_pes_14_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_17_clock = clock;
  assign local_pes_14_17_reset = reset;
  assign local_pes_14_17_io_in_q = local_pes_14_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_17_io_in_sum = local_pes_14_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_17_io_in_sum_exp = local_pes_14_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_17_io_in_kv = local_pes_13_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_17_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_17_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_17_io_in_stage = local_pes_14_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_18_clock = clock;
  assign local_pes_14_18_reset = reset;
  assign local_pes_14_18_io_in_q = local_pes_14_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_18_io_in_sum = local_pes_14_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_18_io_in_sum_exp = local_pes_14_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_18_io_in_kv = local_pes_13_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_18_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_18_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_18_io_in_stage = local_pes_14_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_19_clock = clock;
  assign local_pes_14_19_reset = reset;
  assign local_pes_14_19_io_in_q = local_pes_14_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_19_io_in_sum = local_pes_14_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_19_io_in_sum_exp = local_pes_14_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_19_io_in_kv = local_pes_13_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_19_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_19_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_19_io_in_stage = local_pes_14_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_20_clock = clock;
  assign local_pes_14_20_reset = reset;
  assign local_pes_14_20_io_in_q = local_pes_14_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_20_io_in_sum = local_pes_14_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_20_io_in_sum_exp = local_pes_14_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_20_io_in_kv = local_pes_13_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_20_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_20_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_20_io_in_stage = local_pes_14_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_21_clock = clock;
  assign local_pes_14_21_reset = reset;
  assign local_pes_14_21_io_in_q = local_pes_14_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_21_io_in_sum = local_pes_14_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_21_io_in_sum_exp = local_pes_14_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_21_io_in_kv = local_pes_13_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_21_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_21_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_21_io_in_stage = local_pes_14_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_22_clock = clock;
  assign local_pes_14_22_reset = reset;
  assign local_pes_14_22_io_in_q = local_pes_14_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_22_io_in_sum = local_pes_14_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_22_io_in_sum_exp = local_pes_14_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_22_io_in_kv = local_pes_13_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_22_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_22_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_22_io_in_stage = local_pes_14_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_23_clock = clock;
  assign local_pes_14_23_reset = reset;
  assign local_pes_14_23_io_in_q = local_pes_14_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_23_io_in_sum = local_pes_14_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_23_io_in_sum_exp = local_pes_14_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_23_io_in_kv = local_pes_13_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_23_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_23_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_23_io_in_stage = local_pes_14_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_24_clock = clock;
  assign local_pes_14_24_reset = reset;
  assign local_pes_14_24_io_in_q = local_pes_14_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_24_io_in_sum = local_pes_14_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_24_io_in_sum_exp = local_pes_14_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_24_io_in_kv = local_pes_13_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_24_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_24_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_24_io_in_stage = local_pes_14_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_25_clock = clock;
  assign local_pes_14_25_reset = reset;
  assign local_pes_14_25_io_in_q = local_pes_14_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_25_io_in_sum = local_pes_14_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_25_io_in_sum_exp = local_pes_14_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_25_io_in_kv = local_pes_13_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_25_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_25_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_25_io_in_stage = local_pes_14_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_26_clock = clock;
  assign local_pes_14_26_reset = reset;
  assign local_pes_14_26_io_in_q = local_pes_14_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_26_io_in_sum = local_pes_14_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_26_io_in_sum_exp = local_pes_14_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_26_io_in_kv = local_pes_13_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_26_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_26_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_26_io_in_stage = local_pes_14_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_27_clock = clock;
  assign local_pes_14_27_reset = reset;
  assign local_pes_14_27_io_in_q = local_pes_14_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_27_io_in_sum = local_pes_14_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_27_io_in_sum_exp = local_pes_14_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_27_io_in_kv = local_pes_13_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_27_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_27_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_27_io_in_stage = local_pes_14_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_28_clock = clock;
  assign local_pes_14_28_reset = reset;
  assign local_pes_14_28_io_in_q = local_pes_14_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_28_io_in_sum = local_pes_14_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_28_io_in_sum_exp = local_pes_14_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_28_io_in_kv = local_pes_13_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_28_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_28_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_28_io_in_stage = local_pes_14_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_29_clock = clock;
  assign local_pes_14_29_reset = reset;
  assign local_pes_14_29_io_in_q = local_pes_14_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_29_io_in_sum = local_pes_14_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_29_io_in_sum_exp = local_pes_14_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_29_io_in_kv = local_pes_13_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_29_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_29_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_29_io_in_stage = local_pes_14_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_30_clock = clock;
  assign local_pes_14_30_reset = reset;
  assign local_pes_14_30_io_in_q = local_pes_14_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_30_io_in_sum = local_pes_14_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_30_io_in_sum_exp = local_pes_14_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_30_io_in_kv = local_pes_13_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_30_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_30_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_30_io_in_stage = local_pes_14_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_14_31_clock = clock;
  assign local_pes_14_31_reset = reset;
  assign local_pes_14_31_io_in_q = local_pes_14_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_14_31_io_in_sum = local_pes_14_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_14_31_io_in_sum_exp = local_pes_14_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_14_31_io_in_kv = local_pes_13_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_14_31_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_14_31_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_14_31_io_in_stage = local_pes_14_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_0_clock = clock;
  assign local_pes_15_0_reset = reset;
  assign local_pes_15_0_io_in_q = io_q_ports_15; // @[PEArray.scala 51:37]
  assign local_pes_15_0_io_in_kv = io_kv_ports_46; // @[PEArray.scala 40:34]
  assign local_pes_15_0_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_0_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_0_io_in_stage = io_stage_ports_15; // @[PEArray.scala 52:41]
  assign local_pes_15_1_clock = clock;
  assign local_pes_15_1_reset = reset;
  assign local_pes_15_1_io_in_q = local_pes_15_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_1_io_in_sum = local_pes_15_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_15_1_io_in_kv = local_pes_14_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_1_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_1_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_1_io_in_stage = local_pes_15_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_2_clock = clock;
  assign local_pes_15_2_reset = reset;
  assign local_pes_15_2_io_in_q = local_pes_15_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_2_io_in_sum = local_pes_15_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_2_io_in_sum_exp = local_pes_15_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_2_io_in_kv = local_pes_14_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_2_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_2_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_2_io_in_stage = local_pes_15_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_3_clock = clock;
  assign local_pes_15_3_reset = reset;
  assign local_pes_15_3_io_in_q = local_pes_15_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_3_io_in_sum = local_pes_15_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_3_io_in_sum_exp = local_pes_15_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_3_io_in_kv = local_pes_14_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_3_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_3_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_3_io_in_stage = local_pes_15_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_4_clock = clock;
  assign local_pes_15_4_reset = reset;
  assign local_pes_15_4_io_in_q = local_pes_15_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_4_io_in_sum = local_pes_15_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_4_io_in_sum_exp = local_pes_15_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_4_io_in_kv = local_pes_14_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_4_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_4_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_4_io_in_stage = local_pes_15_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_5_clock = clock;
  assign local_pes_15_5_reset = reset;
  assign local_pes_15_5_io_in_q = local_pes_15_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_5_io_in_sum = local_pes_15_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_5_io_in_sum_exp = local_pes_15_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_5_io_in_kv = local_pes_14_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_5_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_5_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_5_io_in_stage = local_pes_15_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_6_clock = clock;
  assign local_pes_15_6_reset = reset;
  assign local_pes_15_6_io_in_q = local_pes_15_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_6_io_in_sum = local_pes_15_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_6_io_in_sum_exp = local_pes_15_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_6_io_in_kv = local_pes_14_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_6_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_6_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_6_io_in_stage = local_pes_15_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_7_clock = clock;
  assign local_pes_15_7_reset = reset;
  assign local_pes_15_7_io_in_q = local_pes_15_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_7_io_in_sum = local_pes_15_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_7_io_in_sum_exp = local_pes_15_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_7_io_in_kv = local_pes_14_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_7_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_7_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_7_io_in_stage = local_pes_15_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_8_clock = clock;
  assign local_pes_15_8_reset = reset;
  assign local_pes_15_8_io_in_q = local_pes_15_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_8_io_in_sum = local_pes_15_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_8_io_in_sum_exp = local_pes_15_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_8_io_in_kv = local_pes_14_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_8_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_8_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_8_io_in_stage = local_pes_15_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_9_clock = clock;
  assign local_pes_15_9_reset = reset;
  assign local_pes_15_9_io_in_q = local_pes_15_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_9_io_in_sum = local_pes_15_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_9_io_in_sum_exp = local_pes_15_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_9_io_in_kv = local_pes_14_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_9_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_9_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_9_io_in_stage = local_pes_15_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_10_clock = clock;
  assign local_pes_15_10_reset = reset;
  assign local_pes_15_10_io_in_q = local_pes_15_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_10_io_in_sum = local_pes_15_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_10_io_in_sum_exp = local_pes_15_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_10_io_in_kv = local_pes_14_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_10_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_10_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_10_io_in_stage = local_pes_15_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_11_clock = clock;
  assign local_pes_15_11_reset = reset;
  assign local_pes_15_11_io_in_q = local_pes_15_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_11_io_in_sum = local_pes_15_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_11_io_in_sum_exp = local_pes_15_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_11_io_in_kv = local_pes_14_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_11_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_11_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_11_io_in_stage = local_pes_15_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_12_clock = clock;
  assign local_pes_15_12_reset = reset;
  assign local_pes_15_12_io_in_q = local_pes_15_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_12_io_in_sum = local_pes_15_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_12_io_in_sum_exp = local_pes_15_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_12_io_in_kv = local_pes_14_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_12_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_12_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_12_io_in_stage = local_pes_15_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_13_clock = clock;
  assign local_pes_15_13_reset = reset;
  assign local_pes_15_13_io_in_q = local_pes_15_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_13_io_in_sum = local_pes_15_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_13_io_in_sum_exp = local_pes_15_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_13_io_in_kv = local_pes_14_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_13_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_13_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_13_io_in_stage = local_pes_15_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_14_clock = clock;
  assign local_pes_15_14_reset = reset;
  assign local_pes_15_14_io_in_q = local_pes_15_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_14_io_in_sum = local_pes_15_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_14_io_in_sum_exp = local_pes_15_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_14_io_in_kv = local_pes_14_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_14_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_14_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_14_io_in_stage = local_pes_15_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_15_clock = clock;
  assign local_pes_15_15_reset = reset;
  assign local_pes_15_15_io_in_q = local_pes_15_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_15_io_in_sum = local_pes_15_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_15_io_in_sum_exp = local_pes_15_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_15_io_in_kv = local_pes_14_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_15_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_15_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_15_io_in_stage = local_pes_15_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_16_clock = clock;
  assign local_pes_15_16_reset = reset;
  assign local_pes_15_16_io_in_q = local_pes_15_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_16_io_in_sum = local_pes_15_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_16_io_in_sum_exp = local_pes_15_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_16_io_in_kv = local_pes_14_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_16_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_16_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_16_io_in_stage = local_pes_15_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_17_clock = clock;
  assign local_pes_15_17_reset = reset;
  assign local_pes_15_17_io_in_q = local_pes_15_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_17_io_in_sum = local_pes_15_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_17_io_in_sum_exp = local_pes_15_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_17_io_in_kv = local_pes_14_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_17_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_17_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_17_io_in_stage = local_pes_15_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_18_clock = clock;
  assign local_pes_15_18_reset = reset;
  assign local_pes_15_18_io_in_q = local_pes_15_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_18_io_in_sum = local_pes_15_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_18_io_in_sum_exp = local_pes_15_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_18_io_in_kv = local_pes_14_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_18_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_18_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_18_io_in_stage = local_pes_15_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_19_clock = clock;
  assign local_pes_15_19_reset = reset;
  assign local_pes_15_19_io_in_q = local_pes_15_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_19_io_in_sum = local_pes_15_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_19_io_in_sum_exp = local_pes_15_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_19_io_in_kv = local_pes_14_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_19_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_19_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_19_io_in_stage = local_pes_15_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_20_clock = clock;
  assign local_pes_15_20_reset = reset;
  assign local_pes_15_20_io_in_q = local_pes_15_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_20_io_in_sum = local_pes_15_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_20_io_in_sum_exp = local_pes_15_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_20_io_in_kv = local_pes_14_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_20_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_20_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_20_io_in_stage = local_pes_15_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_21_clock = clock;
  assign local_pes_15_21_reset = reset;
  assign local_pes_15_21_io_in_q = local_pes_15_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_21_io_in_sum = local_pes_15_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_21_io_in_sum_exp = local_pes_15_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_21_io_in_kv = local_pes_14_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_21_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_21_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_21_io_in_stage = local_pes_15_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_22_clock = clock;
  assign local_pes_15_22_reset = reset;
  assign local_pes_15_22_io_in_q = local_pes_15_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_22_io_in_sum = local_pes_15_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_22_io_in_sum_exp = local_pes_15_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_22_io_in_kv = local_pes_14_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_22_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_22_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_22_io_in_stage = local_pes_15_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_23_clock = clock;
  assign local_pes_15_23_reset = reset;
  assign local_pes_15_23_io_in_q = local_pes_15_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_23_io_in_sum = local_pes_15_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_23_io_in_sum_exp = local_pes_15_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_23_io_in_kv = local_pes_14_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_23_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_23_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_23_io_in_stage = local_pes_15_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_24_clock = clock;
  assign local_pes_15_24_reset = reset;
  assign local_pes_15_24_io_in_q = local_pes_15_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_24_io_in_sum = local_pes_15_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_24_io_in_sum_exp = local_pes_15_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_24_io_in_kv = local_pes_14_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_24_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_24_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_24_io_in_stage = local_pes_15_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_25_clock = clock;
  assign local_pes_15_25_reset = reset;
  assign local_pes_15_25_io_in_q = local_pes_15_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_25_io_in_sum = local_pes_15_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_25_io_in_sum_exp = local_pes_15_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_25_io_in_kv = local_pes_14_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_25_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_25_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_25_io_in_stage = local_pes_15_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_26_clock = clock;
  assign local_pes_15_26_reset = reset;
  assign local_pes_15_26_io_in_q = local_pes_15_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_26_io_in_sum = local_pes_15_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_26_io_in_sum_exp = local_pes_15_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_26_io_in_kv = local_pes_14_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_26_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_26_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_26_io_in_stage = local_pes_15_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_27_clock = clock;
  assign local_pes_15_27_reset = reset;
  assign local_pes_15_27_io_in_q = local_pes_15_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_27_io_in_sum = local_pes_15_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_27_io_in_sum_exp = local_pes_15_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_27_io_in_kv = local_pes_14_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_27_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_27_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_27_io_in_stage = local_pes_15_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_28_clock = clock;
  assign local_pes_15_28_reset = reset;
  assign local_pes_15_28_io_in_q = local_pes_15_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_28_io_in_sum = local_pes_15_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_28_io_in_sum_exp = local_pes_15_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_28_io_in_kv = local_pes_14_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_28_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_28_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_28_io_in_stage = local_pes_15_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_29_clock = clock;
  assign local_pes_15_29_reset = reset;
  assign local_pes_15_29_io_in_q = local_pes_15_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_29_io_in_sum = local_pes_15_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_29_io_in_sum_exp = local_pes_15_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_29_io_in_kv = local_pes_14_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_29_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_29_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_29_io_in_stage = local_pes_15_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_30_clock = clock;
  assign local_pes_15_30_reset = reset;
  assign local_pes_15_30_io_in_q = local_pes_15_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_30_io_in_sum = local_pes_15_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_30_io_in_sum_exp = local_pes_15_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_30_io_in_kv = local_pes_14_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_30_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_30_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_30_io_in_stage = local_pes_15_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_15_31_clock = clock;
  assign local_pes_15_31_reset = reset;
  assign local_pes_15_31_io_in_q = local_pes_15_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_15_31_io_in_sum = local_pes_15_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_15_31_io_in_sum_exp = local_pes_15_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_15_31_io_in_kv = local_pes_14_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_15_31_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_15_31_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_15_31_io_in_stage = local_pes_15_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_0_clock = clock;
  assign local_pes_16_0_reset = reset;
  assign local_pes_16_0_io_in_q = io_q_ports_16; // @[PEArray.scala 51:37]
  assign local_pes_16_0_io_in_kv = io_kv_ports_47; // @[PEArray.scala 40:34]
  assign local_pes_16_0_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_0_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_0_io_in_stage = io_stage_ports_16; // @[PEArray.scala 52:41]
  assign local_pes_16_1_clock = clock;
  assign local_pes_16_1_reset = reset;
  assign local_pes_16_1_io_in_q = local_pes_16_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_1_io_in_sum = local_pes_16_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_16_1_io_in_kv = local_pes_15_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_1_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_1_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_1_io_in_stage = local_pes_16_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_2_clock = clock;
  assign local_pes_16_2_reset = reset;
  assign local_pes_16_2_io_in_q = local_pes_16_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_2_io_in_sum = local_pes_16_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_2_io_in_sum_exp = local_pes_16_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_2_io_in_kv = local_pes_15_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_2_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_2_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_2_io_in_stage = local_pes_16_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_3_clock = clock;
  assign local_pes_16_3_reset = reset;
  assign local_pes_16_3_io_in_q = local_pes_16_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_3_io_in_sum = local_pes_16_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_3_io_in_sum_exp = local_pes_16_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_3_io_in_kv = local_pes_15_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_3_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_3_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_3_io_in_stage = local_pes_16_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_4_clock = clock;
  assign local_pes_16_4_reset = reset;
  assign local_pes_16_4_io_in_q = local_pes_16_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_4_io_in_sum = local_pes_16_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_4_io_in_sum_exp = local_pes_16_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_4_io_in_kv = local_pes_15_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_4_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_4_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_4_io_in_stage = local_pes_16_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_5_clock = clock;
  assign local_pes_16_5_reset = reset;
  assign local_pes_16_5_io_in_q = local_pes_16_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_5_io_in_sum = local_pes_16_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_5_io_in_sum_exp = local_pes_16_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_5_io_in_kv = local_pes_15_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_5_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_5_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_5_io_in_stage = local_pes_16_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_6_clock = clock;
  assign local_pes_16_6_reset = reset;
  assign local_pes_16_6_io_in_q = local_pes_16_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_6_io_in_sum = local_pes_16_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_6_io_in_sum_exp = local_pes_16_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_6_io_in_kv = local_pes_15_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_6_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_6_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_6_io_in_stage = local_pes_16_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_7_clock = clock;
  assign local_pes_16_7_reset = reset;
  assign local_pes_16_7_io_in_q = local_pes_16_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_7_io_in_sum = local_pes_16_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_7_io_in_sum_exp = local_pes_16_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_7_io_in_kv = local_pes_15_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_7_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_7_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_7_io_in_stage = local_pes_16_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_8_clock = clock;
  assign local_pes_16_8_reset = reset;
  assign local_pes_16_8_io_in_q = local_pes_16_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_8_io_in_sum = local_pes_16_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_8_io_in_sum_exp = local_pes_16_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_8_io_in_kv = local_pes_15_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_8_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_8_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_8_io_in_stage = local_pes_16_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_9_clock = clock;
  assign local_pes_16_9_reset = reset;
  assign local_pes_16_9_io_in_q = local_pes_16_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_9_io_in_sum = local_pes_16_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_9_io_in_sum_exp = local_pes_16_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_9_io_in_kv = local_pes_15_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_9_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_9_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_9_io_in_stage = local_pes_16_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_10_clock = clock;
  assign local_pes_16_10_reset = reset;
  assign local_pes_16_10_io_in_q = local_pes_16_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_10_io_in_sum = local_pes_16_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_10_io_in_sum_exp = local_pes_16_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_10_io_in_kv = local_pes_15_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_10_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_10_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_10_io_in_stage = local_pes_16_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_11_clock = clock;
  assign local_pes_16_11_reset = reset;
  assign local_pes_16_11_io_in_q = local_pes_16_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_11_io_in_sum = local_pes_16_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_11_io_in_sum_exp = local_pes_16_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_11_io_in_kv = local_pes_15_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_11_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_11_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_11_io_in_stage = local_pes_16_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_12_clock = clock;
  assign local_pes_16_12_reset = reset;
  assign local_pes_16_12_io_in_q = local_pes_16_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_12_io_in_sum = local_pes_16_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_12_io_in_sum_exp = local_pes_16_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_12_io_in_kv = local_pes_15_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_12_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_12_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_12_io_in_stage = local_pes_16_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_13_clock = clock;
  assign local_pes_16_13_reset = reset;
  assign local_pes_16_13_io_in_q = local_pes_16_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_13_io_in_sum = local_pes_16_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_13_io_in_sum_exp = local_pes_16_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_13_io_in_kv = local_pes_15_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_13_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_13_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_13_io_in_stage = local_pes_16_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_14_clock = clock;
  assign local_pes_16_14_reset = reset;
  assign local_pes_16_14_io_in_q = local_pes_16_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_14_io_in_sum = local_pes_16_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_14_io_in_sum_exp = local_pes_16_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_14_io_in_kv = local_pes_15_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_14_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_14_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_14_io_in_stage = local_pes_16_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_15_clock = clock;
  assign local_pes_16_15_reset = reset;
  assign local_pes_16_15_io_in_q = local_pes_16_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_15_io_in_sum = local_pes_16_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_15_io_in_sum_exp = local_pes_16_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_15_io_in_kv = local_pes_15_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_15_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_15_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_15_io_in_stage = local_pes_16_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_16_clock = clock;
  assign local_pes_16_16_reset = reset;
  assign local_pes_16_16_io_in_q = local_pes_16_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_16_io_in_sum = local_pes_16_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_16_io_in_sum_exp = local_pes_16_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_16_io_in_kv = local_pes_15_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_16_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_16_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_16_io_in_stage = local_pes_16_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_17_clock = clock;
  assign local_pes_16_17_reset = reset;
  assign local_pes_16_17_io_in_q = local_pes_16_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_17_io_in_sum = local_pes_16_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_17_io_in_sum_exp = local_pes_16_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_17_io_in_kv = local_pes_15_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_17_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_17_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_17_io_in_stage = local_pes_16_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_18_clock = clock;
  assign local_pes_16_18_reset = reset;
  assign local_pes_16_18_io_in_q = local_pes_16_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_18_io_in_sum = local_pes_16_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_18_io_in_sum_exp = local_pes_16_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_18_io_in_kv = local_pes_15_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_18_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_18_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_18_io_in_stage = local_pes_16_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_19_clock = clock;
  assign local_pes_16_19_reset = reset;
  assign local_pes_16_19_io_in_q = local_pes_16_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_19_io_in_sum = local_pes_16_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_19_io_in_sum_exp = local_pes_16_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_19_io_in_kv = local_pes_15_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_19_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_19_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_19_io_in_stage = local_pes_16_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_20_clock = clock;
  assign local_pes_16_20_reset = reset;
  assign local_pes_16_20_io_in_q = local_pes_16_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_20_io_in_sum = local_pes_16_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_20_io_in_sum_exp = local_pes_16_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_20_io_in_kv = local_pes_15_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_20_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_20_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_20_io_in_stage = local_pes_16_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_21_clock = clock;
  assign local_pes_16_21_reset = reset;
  assign local_pes_16_21_io_in_q = local_pes_16_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_21_io_in_sum = local_pes_16_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_21_io_in_sum_exp = local_pes_16_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_21_io_in_kv = local_pes_15_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_21_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_21_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_21_io_in_stage = local_pes_16_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_22_clock = clock;
  assign local_pes_16_22_reset = reset;
  assign local_pes_16_22_io_in_q = local_pes_16_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_22_io_in_sum = local_pes_16_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_22_io_in_sum_exp = local_pes_16_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_22_io_in_kv = local_pes_15_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_22_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_22_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_22_io_in_stage = local_pes_16_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_23_clock = clock;
  assign local_pes_16_23_reset = reset;
  assign local_pes_16_23_io_in_q = local_pes_16_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_23_io_in_sum = local_pes_16_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_23_io_in_sum_exp = local_pes_16_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_23_io_in_kv = local_pes_15_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_23_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_23_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_23_io_in_stage = local_pes_16_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_24_clock = clock;
  assign local_pes_16_24_reset = reset;
  assign local_pes_16_24_io_in_q = local_pes_16_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_24_io_in_sum = local_pes_16_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_24_io_in_sum_exp = local_pes_16_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_24_io_in_kv = local_pes_15_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_24_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_24_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_24_io_in_stage = local_pes_16_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_25_clock = clock;
  assign local_pes_16_25_reset = reset;
  assign local_pes_16_25_io_in_q = local_pes_16_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_25_io_in_sum = local_pes_16_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_25_io_in_sum_exp = local_pes_16_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_25_io_in_kv = local_pes_15_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_25_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_25_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_25_io_in_stage = local_pes_16_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_26_clock = clock;
  assign local_pes_16_26_reset = reset;
  assign local_pes_16_26_io_in_q = local_pes_16_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_26_io_in_sum = local_pes_16_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_26_io_in_sum_exp = local_pes_16_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_26_io_in_kv = local_pes_15_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_26_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_26_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_26_io_in_stage = local_pes_16_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_27_clock = clock;
  assign local_pes_16_27_reset = reset;
  assign local_pes_16_27_io_in_q = local_pes_16_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_27_io_in_sum = local_pes_16_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_27_io_in_sum_exp = local_pes_16_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_27_io_in_kv = local_pes_15_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_27_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_27_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_27_io_in_stage = local_pes_16_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_28_clock = clock;
  assign local_pes_16_28_reset = reset;
  assign local_pes_16_28_io_in_q = local_pes_16_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_28_io_in_sum = local_pes_16_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_28_io_in_sum_exp = local_pes_16_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_28_io_in_kv = local_pes_15_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_28_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_28_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_28_io_in_stage = local_pes_16_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_29_clock = clock;
  assign local_pes_16_29_reset = reset;
  assign local_pes_16_29_io_in_q = local_pes_16_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_29_io_in_sum = local_pes_16_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_29_io_in_sum_exp = local_pes_16_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_29_io_in_kv = local_pes_15_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_29_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_29_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_29_io_in_stage = local_pes_16_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_30_clock = clock;
  assign local_pes_16_30_reset = reset;
  assign local_pes_16_30_io_in_q = local_pes_16_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_30_io_in_sum = local_pes_16_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_30_io_in_sum_exp = local_pes_16_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_30_io_in_kv = local_pes_15_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_30_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_30_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_30_io_in_stage = local_pes_16_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_16_31_clock = clock;
  assign local_pes_16_31_reset = reset;
  assign local_pes_16_31_io_in_q = local_pes_16_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_16_31_io_in_sum = local_pes_16_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_16_31_io_in_sum_exp = local_pes_16_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_16_31_io_in_kv = local_pes_15_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_16_31_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_16_31_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_16_31_io_in_stage = local_pes_16_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_0_clock = clock;
  assign local_pes_17_0_reset = reset;
  assign local_pes_17_0_io_in_q = io_q_ports_17; // @[PEArray.scala 51:37]
  assign local_pes_17_0_io_in_kv = io_kv_ports_48; // @[PEArray.scala 40:34]
  assign local_pes_17_0_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_0_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_0_io_in_stage = io_stage_ports_17; // @[PEArray.scala 52:41]
  assign local_pes_17_1_clock = clock;
  assign local_pes_17_1_reset = reset;
  assign local_pes_17_1_io_in_q = local_pes_17_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_1_io_in_sum = local_pes_17_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_17_1_io_in_kv = local_pes_16_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_1_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_1_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_1_io_in_stage = local_pes_17_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_2_clock = clock;
  assign local_pes_17_2_reset = reset;
  assign local_pes_17_2_io_in_q = local_pes_17_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_2_io_in_sum = local_pes_17_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_2_io_in_sum_exp = local_pes_17_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_2_io_in_kv = local_pes_16_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_2_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_2_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_2_io_in_stage = local_pes_17_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_3_clock = clock;
  assign local_pes_17_3_reset = reset;
  assign local_pes_17_3_io_in_q = local_pes_17_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_3_io_in_sum = local_pes_17_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_3_io_in_sum_exp = local_pes_17_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_3_io_in_kv = local_pes_16_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_3_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_3_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_3_io_in_stage = local_pes_17_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_4_clock = clock;
  assign local_pes_17_4_reset = reset;
  assign local_pes_17_4_io_in_q = local_pes_17_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_4_io_in_sum = local_pes_17_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_4_io_in_sum_exp = local_pes_17_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_4_io_in_kv = local_pes_16_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_4_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_4_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_4_io_in_stage = local_pes_17_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_5_clock = clock;
  assign local_pes_17_5_reset = reset;
  assign local_pes_17_5_io_in_q = local_pes_17_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_5_io_in_sum = local_pes_17_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_5_io_in_sum_exp = local_pes_17_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_5_io_in_kv = local_pes_16_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_5_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_5_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_5_io_in_stage = local_pes_17_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_6_clock = clock;
  assign local_pes_17_6_reset = reset;
  assign local_pes_17_6_io_in_q = local_pes_17_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_6_io_in_sum = local_pes_17_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_6_io_in_sum_exp = local_pes_17_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_6_io_in_kv = local_pes_16_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_6_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_6_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_6_io_in_stage = local_pes_17_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_7_clock = clock;
  assign local_pes_17_7_reset = reset;
  assign local_pes_17_7_io_in_q = local_pes_17_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_7_io_in_sum = local_pes_17_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_7_io_in_sum_exp = local_pes_17_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_7_io_in_kv = local_pes_16_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_7_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_7_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_7_io_in_stage = local_pes_17_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_8_clock = clock;
  assign local_pes_17_8_reset = reset;
  assign local_pes_17_8_io_in_q = local_pes_17_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_8_io_in_sum = local_pes_17_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_8_io_in_sum_exp = local_pes_17_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_8_io_in_kv = local_pes_16_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_8_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_8_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_8_io_in_stage = local_pes_17_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_9_clock = clock;
  assign local_pes_17_9_reset = reset;
  assign local_pes_17_9_io_in_q = local_pes_17_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_9_io_in_sum = local_pes_17_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_9_io_in_sum_exp = local_pes_17_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_9_io_in_kv = local_pes_16_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_9_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_9_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_9_io_in_stage = local_pes_17_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_10_clock = clock;
  assign local_pes_17_10_reset = reset;
  assign local_pes_17_10_io_in_q = local_pes_17_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_10_io_in_sum = local_pes_17_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_10_io_in_sum_exp = local_pes_17_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_10_io_in_kv = local_pes_16_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_10_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_10_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_10_io_in_stage = local_pes_17_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_11_clock = clock;
  assign local_pes_17_11_reset = reset;
  assign local_pes_17_11_io_in_q = local_pes_17_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_11_io_in_sum = local_pes_17_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_11_io_in_sum_exp = local_pes_17_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_11_io_in_kv = local_pes_16_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_11_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_11_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_11_io_in_stage = local_pes_17_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_12_clock = clock;
  assign local_pes_17_12_reset = reset;
  assign local_pes_17_12_io_in_q = local_pes_17_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_12_io_in_sum = local_pes_17_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_12_io_in_sum_exp = local_pes_17_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_12_io_in_kv = local_pes_16_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_12_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_12_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_12_io_in_stage = local_pes_17_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_13_clock = clock;
  assign local_pes_17_13_reset = reset;
  assign local_pes_17_13_io_in_q = local_pes_17_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_13_io_in_sum = local_pes_17_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_13_io_in_sum_exp = local_pes_17_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_13_io_in_kv = local_pes_16_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_13_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_13_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_13_io_in_stage = local_pes_17_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_14_clock = clock;
  assign local_pes_17_14_reset = reset;
  assign local_pes_17_14_io_in_q = local_pes_17_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_14_io_in_sum = local_pes_17_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_14_io_in_sum_exp = local_pes_17_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_14_io_in_kv = local_pes_16_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_14_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_14_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_14_io_in_stage = local_pes_17_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_15_clock = clock;
  assign local_pes_17_15_reset = reset;
  assign local_pes_17_15_io_in_q = local_pes_17_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_15_io_in_sum = local_pes_17_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_15_io_in_sum_exp = local_pes_17_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_15_io_in_kv = local_pes_16_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_15_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_15_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_15_io_in_stage = local_pes_17_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_16_clock = clock;
  assign local_pes_17_16_reset = reset;
  assign local_pes_17_16_io_in_q = local_pes_17_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_16_io_in_sum = local_pes_17_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_16_io_in_sum_exp = local_pes_17_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_16_io_in_kv = local_pes_16_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_16_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_16_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_16_io_in_stage = local_pes_17_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_17_clock = clock;
  assign local_pes_17_17_reset = reset;
  assign local_pes_17_17_io_in_q = local_pes_17_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_17_io_in_sum = local_pes_17_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_17_io_in_sum_exp = local_pes_17_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_17_io_in_kv = local_pes_16_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_17_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_17_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_17_io_in_stage = local_pes_17_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_18_clock = clock;
  assign local_pes_17_18_reset = reset;
  assign local_pes_17_18_io_in_q = local_pes_17_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_18_io_in_sum = local_pes_17_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_18_io_in_sum_exp = local_pes_17_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_18_io_in_kv = local_pes_16_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_18_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_18_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_18_io_in_stage = local_pes_17_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_19_clock = clock;
  assign local_pes_17_19_reset = reset;
  assign local_pes_17_19_io_in_q = local_pes_17_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_19_io_in_sum = local_pes_17_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_19_io_in_sum_exp = local_pes_17_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_19_io_in_kv = local_pes_16_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_19_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_19_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_19_io_in_stage = local_pes_17_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_20_clock = clock;
  assign local_pes_17_20_reset = reset;
  assign local_pes_17_20_io_in_q = local_pes_17_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_20_io_in_sum = local_pes_17_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_20_io_in_sum_exp = local_pes_17_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_20_io_in_kv = local_pes_16_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_20_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_20_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_20_io_in_stage = local_pes_17_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_21_clock = clock;
  assign local_pes_17_21_reset = reset;
  assign local_pes_17_21_io_in_q = local_pes_17_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_21_io_in_sum = local_pes_17_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_21_io_in_sum_exp = local_pes_17_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_21_io_in_kv = local_pes_16_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_21_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_21_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_21_io_in_stage = local_pes_17_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_22_clock = clock;
  assign local_pes_17_22_reset = reset;
  assign local_pes_17_22_io_in_q = local_pes_17_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_22_io_in_sum = local_pes_17_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_22_io_in_sum_exp = local_pes_17_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_22_io_in_kv = local_pes_16_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_22_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_22_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_22_io_in_stage = local_pes_17_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_23_clock = clock;
  assign local_pes_17_23_reset = reset;
  assign local_pes_17_23_io_in_q = local_pes_17_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_23_io_in_sum = local_pes_17_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_23_io_in_sum_exp = local_pes_17_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_23_io_in_kv = local_pes_16_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_23_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_23_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_23_io_in_stage = local_pes_17_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_24_clock = clock;
  assign local_pes_17_24_reset = reset;
  assign local_pes_17_24_io_in_q = local_pes_17_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_24_io_in_sum = local_pes_17_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_24_io_in_sum_exp = local_pes_17_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_24_io_in_kv = local_pes_16_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_24_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_24_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_24_io_in_stage = local_pes_17_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_25_clock = clock;
  assign local_pes_17_25_reset = reset;
  assign local_pes_17_25_io_in_q = local_pes_17_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_25_io_in_sum = local_pes_17_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_25_io_in_sum_exp = local_pes_17_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_25_io_in_kv = local_pes_16_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_25_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_25_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_25_io_in_stage = local_pes_17_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_26_clock = clock;
  assign local_pes_17_26_reset = reset;
  assign local_pes_17_26_io_in_q = local_pes_17_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_26_io_in_sum = local_pes_17_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_26_io_in_sum_exp = local_pes_17_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_26_io_in_kv = local_pes_16_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_26_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_26_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_26_io_in_stage = local_pes_17_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_27_clock = clock;
  assign local_pes_17_27_reset = reset;
  assign local_pes_17_27_io_in_q = local_pes_17_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_27_io_in_sum = local_pes_17_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_27_io_in_sum_exp = local_pes_17_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_27_io_in_kv = local_pes_16_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_27_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_27_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_27_io_in_stage = local_pes_17_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_28_clock = clock;
  assign local_pes_17_28_reset = reset;
  assign local_pes_17_28_io_in_q = local_pes_17_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_28_io_in_sum = local_pes_17_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_28_io_in_sum_exp = local_pes_17_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_28_io_in_kv = local_pes_16_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_28_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_28_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_28_io_in_stage = local_pes_17_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_29_clock = clock;
  assign local_pes_17_29_reset = reset;
  assign local_pes_17_29_io_in_q = local_pes_17_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_29_io_in_sum = local_pes_17_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_29_io_in_sum_exp = local_pes_17_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_29_io_in_kv = local_pes_16_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_29_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_29_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_29_io_in_stage = local_pes_17_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_30_clock = clock;
  assign local_pes_17_30_reset = reset;
  assign local_pes_17_30_io_in_q = local_pes_17_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_30_io_in_sum = local_pes_17_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_30_io_in_sum_exp = local_pes_17_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_30_io_in_kv = local_pes_16_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_30_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_30_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_30_io_in_stage = local_pes_17_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_17_31_clock = clock;
  assign local_pes_17_31_reset = reset;
  assign local_pes_17_31_io_in_q = local_pes_17_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_17_31_io_in_sum = local_pes_17_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_17_31_io_in_sum_exp = local_pes_17_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_17_31_io_in_kv = local_pes_16_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_17_31_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_17_31_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_17_31_io_in_stage = local_pes_17_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_0_clock = clock;
  assign local_pes_18_0_reset = reset;
  assign local_pes_18_0_io_in_q = io_q_ports_18; // @[PEArray.scala 51:37]
  assign local_pes_18_0_io_in_kv = io_kv_ports_49; // @[PEArray.scala 40:34]
  assign local_pes_18_0_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_0_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_0_io_in_stage = io_stage_ports_18; // @[PEArray.scala 52:41]
  assign local_pes_18_1_clock = clock;
  assign local_pes_18_1_reset = reset;
  assign local_pes_18_1_io_in_q = local_pes_18_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_1_io_in_sum = local_pes_18_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_18_1_io_in_kv = local_pes_17_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_1_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_1_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_1_io_in_stage = local_pes_18_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_2_clock = clock;
  assign local_pes_18_2_reset = reset;
  assign local_pes_18_2_io_in_q = local_pes_18_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_2_io_in_sum = local_pes_18_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_2_io_in_sum_exp = local_pes_18_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_2_io_in_kv = local_pes_17_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_2_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_2_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_2_io_in_stage = local_pes_18_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_3_clock = clock;
  assign local_pes_18_3_reset = reset;
  assign local_pes_18_3_io_in_q = local_pes_18_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_3_io_in_sum = local_pes_18_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_3_io_in_sum_exp = local_pes_18_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_3_io_in_kv = local_pes_17_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_3_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_3_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_3_io_in_stage = local_pes_18_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_4_clock = clock;
  assign local_pes_18_4_reset = reset;
  assign local_pes_18_4_io_in_q = local_pes_18_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_4_io_in_sum = local_pes_18_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_4_io_in_sum_exp = local_pes_18_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_4_io_in_kv = local_pes_17_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_4_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_4_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_4_io_in_stage = local_pes_18_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_5_clock = clock;
  assign local_pes_18_5_reset = reset;
  assign local_pes_18_5_io_in_q = local_pes_18_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_5_io_in_sum = local_pes_18_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_5_io_in_sum_exp = local_pes_18_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_5_io_in_kv = local_pes_17_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_5_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_5_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_5_io_in_stage = local_pes_18_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_6_clock = clock;
  assign local_pes_18_6_reset = reset;
  assign local_pes_18_6_io_in_q = local_pes_18_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_6_io_in_sum = local_pes_18_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_6_io_in_sum_exp = local_pes_18_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_6_io_in_kv = local_pes_17_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_6_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_6_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_6_io_in_stage = local_pes_18_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_7_clock = clock;
  assign local_pes_18_7_reset = reset;
  assign local_pes_18_7_io_in_q = local_pes_18_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_7_io_in_sum = local_pes_18_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_7_io_in_sum_exp = local_pes_18_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_7_io_in_kv = local_pes_17_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_7_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_7_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_7_io_in_stage = local_pes_18_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_8_clock = clock;
  assign local_pes_18_8_reset = reset;
  assign local_pes_18_8_io_in_q = local_pes_18_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_8_io_in_sum = local_pes_18_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_8_io_in_sum_exp = local_pes_18_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_8_io_in_kv = local_pes_17_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_8_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_8_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_8_io_in_stage = local_pes_18_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_9_clock = clock;
  assign local_pes_18_9_reset = reset;
  assign local_pes_18_9_io_in_q = local_pes_18_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_9_io_in_sum = local_pes_18_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_9_io_in_sum_exp = local_pes_18_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_9_io_in_kv = local_pes_17_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_9_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_9_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_9_io_in_stage = local_pes_18_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_10_clock = clock;
  assign local_pes_18_10_reset = reset;
  assign local_pes_18_10_io_in_q = local_pes_18_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_10_io_in_sum = local_pes_18_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_10_io_in_sum_exp = local_pes_18_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_10_io_in_kv = local_pes_17_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_10_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_10_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_10_io_in_stage = local_pes_18_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_11_clock = clock;
  assign local_pes_18_11_reset = reset;
  assign local_pes_18_11_io_in_q = local_pes_18_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_11_io_in_sum = local_pes_18_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_11_io_in_sum_exp = local_pes_18_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_11_io_in_kv = local_pes_17_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_11_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_11_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_11_io_in_stage = local_pes_18_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_12_clock = clock;
  assign local_pes_18_12_reset = reset;
  assign local_pes_18_12_io_in_q = local_pes_18_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_12_io_in_sum = local_pes_18_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_12_io_in_sum_exp = local_pes_18_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_12_io_in_kv = local_pes_17_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_12_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_12_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_12_io_in_stage = local_pes_18_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_13_clock = clock;
  assign local_pes_18_13_reset = reset;
  assign local_pes_18_13_io_in_q = local_pes_18_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_13_io_in_sum = local_pes_18_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_13_io_in_sum_exp = local_pes_18_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_13_io_in_kv = local_pes_17_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_13_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_13_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_13_io_in_stage = local_pes_18_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_14_clock = clock;
  assign local_pes_18_14_reset = reset;
  assign local_pes_18_14_io_in_q = local_pes_18_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_14_io_in_sum = local_pes_18_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_14_io_in_sum_exp = local_pes_18_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_14_io_in_kv = local_pes_17_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_14_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_14_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_14_io_in_stage = local_pes_18_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_15_clock = clock;
  assign local_pes_18_15_reset = reset;
  assign local_pes_18_15_io_in_q = local_pes_18_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_15_io_in_sum = local_pes_18_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_15_io_in_sum_exp = local_pes_18_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_15_io_in_kv = local_pes_17_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_15_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_15_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_15_io_in_stage = local_pes_18_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_16_clock = clock;
  assign local_pes_18_16_reset = reset;
  assign local_pes_18_16_io_in_q = local_pes_18_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_16_io_in_sum = local_pes_18_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_16_io_in_sum_exp = local_pes_18_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_16_io_in_kv = local_pes_17_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_16_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_16_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_16_io_in_stage = local_pes_18_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_17_clock = clock;
  assign local_pes_18_17_reset = reset;
  assign local_pes_18_17_io_in_q = local_pes_18_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_17_io_in_sum = local_pes_18_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_17_io_in_sum_exp = local_pes_18_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_17_io_in_kv = local_pes_17_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_17_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_17_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_17_io_in_stage = local_pes_18_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_18_clock = clock;
  assign local_pes_18_18_reset = reset;
  assign local_pes_18_18_io_in_q = local_pes_18_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_18_io_in_sum = local_pes_18_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_18_io_in_sum_exp = local_pes_18_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_18_io_in_kv = local_pes_17_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_18_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_18_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_18_io_in_stage = local_pes_18_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_19_clock = clock;
  assign local_pes_18_19_reset = reset;
  assign local_pes_18_19_io_in_q = local_pes_18_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_19_io_in_sum = local_pes_18_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_19_io_in_sum_exp = local_pes_18_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_19_io_in_kv = local_pes_17_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_19_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_19_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_19_io_in_stage = local_pes_18_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_20_clock = clock;
  assign local_pes_18_20_reset = reset;
  assign local_pes_18_20_io_in_q = local_pes_18_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_20_io_in_sum = local_pes_18_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_20_io_in_sum_exp = local_pes_18_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_20_io_in_kv = local_pes_17_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_20_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_20_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_20_io_in_stage = local_pes_18_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_21_clock = clock;
  assign local_pes_18_21_reset = reset;
  assign local_pes_18_21_io_in_q = local_pes_18_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_21_io_in_sum = local_pes_18_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_21_io_in_sum_exp = local_pes_18_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_21_io_in_kv = local_pes_17_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_21_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_21_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_21_io_in_stage = local_pes_18_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_22_clock = clock;
  assign local_pes_18_22_reset = reset;
  assign local_pes_18_22_io_in_q = local_pes_18_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_22_io_in_sum = local_pes_18_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_22_io_in_sum_exp = local_pes_18_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_22_io_in_kv = local_pes_17_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_22_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_22_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_22_io_in_stage = local_pes_18_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_23_clock = clock;
  assign local_pes_18_23_reset = reset;
  assign local_pes_18_23_io_in_q = local_pes_18_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_23_io_in_sum = local_pes_18_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_23_io_in_sum_exp = local_pes_18_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_23_io_in_kv = local_pes_17_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_23_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_23_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_23_io_in_stage = local_pes_18_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_24_clock = clock;
  assign local_pes_18_24_reset = reset;
  assign local_pes_18_24_io_in_q = local_pes_18_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_24_io_in_sum = local_pes_18_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_24_io_in_sum_exp = local_pes_18_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_24_io_in_kv = local_pes_17_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_24_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_24_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_24_io_in_stage = local_pes_18_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_25_clock = clock;
  assign local_pes_18_25_reset = reset;
  assign local_pes_18_25_io_in_q = local_pes_18_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_25_io_in_sum = local_pes_18_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_25_io_in_sum_exp = local_pes_18_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_25_io_in_kv = local_pes_17_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_25_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_25_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_25_io_in_stage = local_pes_18_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_26_clock = clock;
  assign local_pes_18_26_reset = reset;
  assign local_pes_18_26_io_in_q = local_pes_18_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_26_io_in_sum = local_pes_18_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_26_io_in_sum_exp = local_pes_18_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_26_io_in_kv = local_pes_17_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_26_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_26_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_26_io_in_stage = local_pes_18_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_27_clock = clock;
  assign local_pes_18_27_reset = reset;
  assign local_pes_18_27_io_in_q = local_pes_18_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_27_io_in_sum = local_pes_18_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_27_io_in_sum_exp = local_pes_18_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_27_io_in_kv = local_pes_17_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_27_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_27_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_27_io_in_stage = local_pes_18_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_28_clock = clock;
  assign local_pes_18_28_reset = reset;
  assign local_pes_18_28_io_in_q = local_pes_18_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_28_io_in_sum = local_pes_18_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_28_io_in_sum_exp = local_pes_18_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_28_io_in_kv = local_pes_17_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_28_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_28_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_28_io_in_stage = local_pes_18_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_29_clock = clock;
  assign local_pes_18_29_reset = reset;
  assign local_pes_18_29_io_in_q = local_pes_18_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_29_io_in_sum = local_pes_18_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_29_io_in_sum_exp = local_pes_18_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_29_io_in_kv = local_pes_17_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_29_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_29_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_29_io_in_stage = local_pes_18_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_30_clock = clock;
  assign local_pes_18_30_reset = reset;
  assign local_pes_18_30_io_in_q = local_pes_18_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_30_io_in_sum = local_pes_18_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_30_io_in_sum_exp = local_pes_18_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_30_io_in_kv = local_pes_17_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_30_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_30_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_30_io_in_stage = local_pes_18_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_18_31_clock = clock;
  assign local_pes_18_31_reset = reset;
  assign local_pes_18_31_io_in_q = local_pes_18_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_18_31_io_in_sum = local_pes_18_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_18_31_io_in_sum_exp = local_pes_18_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_18_31_io_in_kv = local_pes_17_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_18_31_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_18_31_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_18_31_io_in_stage = local_pes_18_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_0_clock = clock;
  assign local_pes_19_0_reset = reset;
  assign local_pes_19_0_io_in_q = io_q_ports_19; // @[PEArray.scala 51:37]
  assign local_pes_19_0_io_in_kv = io_kv_ports_50; // @[PEArray.scala 40:34]
  assign local_pes_19_0_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_0_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_0_io_in_stage = io_stage_ports_19; // @[PEArray.scala 52:41]
  assign local_pes_19_1_clock = clock;
  assign local_pes_19_1_reset = reset;
  assign local_pes_19_1_io_in_q = local_pes_19_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_1_io_in_sum = local_pes_19_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_19_1_io_in_kv = local_pes_18_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_1_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_1_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_1_io_in_stage = local_pes_19_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_2_clock = clock;
  assign local_pes_19_2_reset = reset;
  assign local_pes_19_2_io_in_q = local_pes_19_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_2_io_in_sum = local_pes_19_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_2_io_in_sum_exp = local_pes_19_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_2_io_in_kv = local_pes_18_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_2_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_2_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_2_io_in_stage = local_pes_19_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_3_clock = clock;
  assign local_pes_19_3_reset = reset;
  assign local_pes_19_3_io_in_q = local_pes_19_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_3_io_in_sum = local_pes_19_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_3_io_in_sum_exp = local_pes_19_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_3_io_in_kv = local_pes_18_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_3_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_3_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_3_io_in_stage = local_pes_19_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_4_clock = clock;
  assign local_pes_19_4_reset = reset;
  assign local_pes_19_4_io_in_q = local_pes_19_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_4_io_in_sum = local_pes_19_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_4_io_in_sum_exp = local_pes_19_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_4_io_in_kv = local_pes_18_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_4_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_4_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_4_io_in_stage = local_pes_19_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_5_clock = clock;
  assign local_pes_19_5_reset = reset;
  assign local_pes_19_5_io_in_q = local_pes_19_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_5_io_in_sum = local_pes_19_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_5_io_in_sum_exp = local_pes_19_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_5_io_in_kv = local_pes_18_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_5_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_5_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_5_io_in_stage = local_pes_19_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_6_clock = clock;
  assign local_pes_19_6_reset = reset;
  assign local_pes_19_6_io_in_q = local_pes_19_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_6_io_in_sum = local_pes_19_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_6_io_in_sum_exp = local_pes_19_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_6_io_in_kv = local_pes_18_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_6_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_6_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_6_io_in_stage = local_pes_19_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_7_clock = clock;
  assign local_pes_19_7_reset = reset;
  assign local_pes_19_7_io_in_q = local_pes_19_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_7_io_in_sum = local_pes_19_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_7_io_in_sum_exp = local_pes_19_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_7_io_in_kv = local_pes_18_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_7_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_7_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_7_io_in_stage = local_pes_19_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_8_clock = clock;
  assign local_pes_19_8_reset = reset;
  assign local_pes_19_8_io_in_q = local_pes_19_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_8_io_in_sum = local_pes_19_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_8_io_in_sum_exp = local_pes_19_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_8_io_in_kv = local_pes_18_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_8_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_8_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_8_io_in_stage = local_pes_19_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_9_clock = clock;
  assign local_pes_19_9_reset = reset;
  assign local_pes_19_9_io_in_q = local_pes_19_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_9_io_in_sum = local_pes_19_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_9_io_in_sum_exp = local_pes_19_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_9_io_in_kv = local_pes_18_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_9_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_9_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_9_io_in_stage = local_pes_19_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_10_clock = clock;
  assign local_pes_19_10_reset = reset;
  assign local_pes_19_10_io_in_q = local_pes_19_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_10_io_in_sum = local_pes_19_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_10_io_in_sum_exp = local_pes_19_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_10_io_in_kv = local_pes_18_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_10_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_10_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_10_io_in_stage = local_pes_19_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_11_clock = clock;
  assign local_pes_19_11_reset = reset;
  assign local_pes_19_11_io_in_q = local_pes_19_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_11_io_in_sum = local_pes_19_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_11_io_in_sum_exp = local_pes_19_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_11_io_in_kv = local_pes_18_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_11_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_11_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_11_io_in_stage = local_pes_19_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_12_clock = clock;
  assign local_pes_19_12_reset = reset;
  assign local_pes_19_12_io_in_q = local_pes_19_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_12_io_in_sum = local_pes_19_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_12_io_in_sum_exp = local_pes_19_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_12_io_in_kv = local_pes_18_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_12_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_12_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_12_io_in_stage = local_pes_19_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_13_clock = clock;
  assign local_pes_19_13_reset = reset;
  assign local_pes_19_13_io_in_q = local_pes_19_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_13_io_in_sum = local_pes_19_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_13_io_in_sum_exp = local_pes_19_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_13_io_in_kv = local_pes_18_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_13_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_13_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_13_io_in_stage = local_pes_19_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_14_clock = clock;
  assign local_pes_19_14_reset = reset;
  assign local_pes_19_14_io_in_q = local_pes_19_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_14_io_in_sum = local_pes_19_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_14_io_in_sum_exp = local_pes_19_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_14_io_in_kv = local_pes_18_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_14_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_14_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_14_io_in_stage = local_pes_19_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_15_clock = clock;
  assign local_pes_19_15_reset = reset;
  assign local_pes_19_15_io_in_q = local_pes_19_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_15_io_in_sum = local_pes_19_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_15_io_in_sum_exp = local_pes_19_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_15_io_in_kv = local_pes_18_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_15_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_15_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_15_io_in_stage = local_pes_19_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_16_clock = clock;
  assign local_pes_19_16_reset = reset;
  assign local_pes_19_16_io_in_q = local_pes_19_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_16_io_in_sum = local_pes_19_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_16_io_in_sum_exp = local_pes_19_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_16_io_in_kv = local_pes_18_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_16_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_16_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_16_io_in_stage = local_pes_19_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_17_clock = clock;
  assign local_pes_19_17_reset = reset;
  assign local_pes_19_17_io_in_q = local_pes_19_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_17_io_in_sum = local_pes_19_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_17_io_in_sum_exp = local_pes_19_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_17_io_in_kv = local_pes_18_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_17_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_17_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_17_io_in_stage = local_pes_19_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_18_clock = clock;
  assign local_pes_19_18_reset = reset;
  assign local_pes_19_18_io_in_q = local_pes_19_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_18_io_in_sum = local_pes_19_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_18_io_in_sum_exp = local_pes_19_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_18_io_in_kv = local_pes_18_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_18_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_18_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_18_io_in_stage = local_pes_19_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_19_clock = clock;
  assign local_pes_19_19_reset = reset;
  assign local_pes_19_19_io_in_q = local_pes_19_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_19_io_in_sum = local_pes_19_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_19_io_in_sum_exp = local_pes_19_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_19_io_in_kv = local_pes_18_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_19_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_19_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_19_io_in_stage = local_pes_19_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_20_clock = clock;
  assign local_pes_19_20_reset = reset;
  assign local_pes_19_20_io_in_q = local_pes_19_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_20_io_in_sum = local_pes_19_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_20_io_in_sum_exp = local_pes_19_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_20_io_in_kv = local_pes_18_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_20_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_20_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_20_io_in_stage = local_pes_19_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_21_clock = clock;
  assign local_pes_19_21_reset = reset;
  assign local_pes_19_21_io_in_q = local_pes_19_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_21_io_in_sum = local_pes_19_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_21_io_in_sum_exp = local_pes_19_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_21_io_in_kv = local_pes_18_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_21_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_21_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_21_io_in_stage = local_pes_19_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_22_clock = clock;
  assign local_pes_19_22_reset = reset;
  assign local_pes_19_22_io_in_q = local_pes_19_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_22_io_in_sum = local_pes_19_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_22_io_in_sum_exp = local_pes_19_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_22_io_in_kv = local_pes_18_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_22_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_22_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_22_io_in_stage = local_pes_19_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_23_clock = clock;
  assign local_pes_19_23_reset = reset;
  assign local_pes_19_23_io_in_q = local_pes_19_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_23_io_in_sum = local_pes_19_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_23_io_in_sum_exp = local_pes_19_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_23_io_in_kv = local_pes_18_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_23_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_23_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_23_io_in_stage = local_pes_19_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_24_clock = clock;
  assign local_pes_19_24_reset = reset;
  assign local_pes_19_24_io_in_q = local_pes_19_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_24_io_in_sum = local_pes_19_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_24_io_in_sum_exp = local_pes_19_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_24_io_in_kv = local_pes_18_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_24_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_24_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_24_io_in_stage = local_pes_19_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_25_clock = clock;
  assign local_pes_19_25_reset = reset;
  assign local_pes_19_25_io_in_q = local_pes_19_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_25_io_in_sum = local_pes_19_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_25_io_in_sum_exp = local_pes_19_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_25_io_in_kv = local_pes_18_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_25_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_25_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_25_io_in_stage = local_pes_19_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_26_clock = clock;
  assign local_pes_19_26_reset = reset;
  assign local_pes_19_26_io_in_q = local_pes_19_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_26_io_in_sum = local_pes_19_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_26_io_in_sum_exp = local_pes_19_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_26_io_in_kv = local_pes_18_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_26_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_26_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_26_io_in_stage = local_pes_19_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_27_clock = clock;
  assign local_pes_19_27_reset = reset;
  assign local_pes_19_27_io_in_q = local_pes_19_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_27_io_in_sum = local_pes_19_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_27_io_in_sum_exp = local_pes_19_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_27_io_in_kv = local_pes_18_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_27_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_27_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_27_io_in_stage = local_pes_19_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_28_clock = clock;
  assign local_pes_19_28_reset = reset;
  assign local_pes_19_28_io_in_q = local_pes_19_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_28_io_in_sum = local_pes_19_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_28_io_in_sum_exp = local_pes_19_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_28_io_in_kv = local_pes_18_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_28_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_28_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_28_io_in_stage = local_pes_19_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_29_clock = clock;
  assign local_pes_19_29_reset = reset;
  assign local_pes_19_29_io_in_q = local_pes_19_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_29_io_in_sum = local_pes_19_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_29_io_in_sum_exp = local_pes_19_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_29_io_in_kv = local_pes_18_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_29_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_29_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_29_io_in_stage = local_pes_19_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_30_clock = clock;
  assign local_pes_19_30_reset = reset;
  assign local_pes_19_30_io_in_q = local_pes_19_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_30_io_in_sum = local_pes_19_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_30_io_in_sum_exp = local_pes_19_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_30_io_in_kv = local_pes_18_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_30_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_30_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_30_io_in_stage = local_pes_19_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_19_31_clock = clock;
  assign local_pes_19_31_reset = reset;
  assign local_pes_19_31_io_in_q = local_pes_19_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_19_31_io_in_sum = local_pes_19_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_19_31_io_in_sum_exp = local_pes_19_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_19_31_io_in_kv = local_pes_18_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_19_31_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_19_31_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_19_31_io_in_stage = local_pes_19_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_0_clock = clock;
  assign local_pes_20_0_reset = reset;
  assign local_pes_20_0_io_in_q = io_q_ports_20; // @[PEArray.scala 51:37]
  assign local_pes_20_0_io_in_kv = io_kv_ports_51; // @[PEArray.scala 40:34]
  assign local_pes_20_0_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_0_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_0_io_in_stage = io_stage_ports_20; // @[PEArray.scala 52:41]
  assign local_pes_20_1_clock = clock;
  assign local_pes_20_1_reset = reset;
  assign local_pes_20_1_io_in_q = local_pes_20_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_1_io_in_sum = local_pes_20_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_20_1_io_in_kv = local_pes_19_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_1_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_1_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_1_io_in_stage = local_pes_20_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_2_clock = clock;
  assign local_pes_20_2_reset = reset;
  assign local_pes_20_2_io_in_q = local_pes_20_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_2_io_in_sum = local_pes_20_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_2_io_in_sum_exp = local_pes_20_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_2_io_in_kv = local_pes_19_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_2_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_2_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_2_io_in_stage = local_pes_20_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_3_clock = clock;
  assign local_pes_20_3_reset = reset;
  assign local_pes_20_3_io_in_q = local_pes_20_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_3_io_in_sum = local_pes_20_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_3_io_in_sum_exp = local_pes_20_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_3_io_in_kv = local_pes_19_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_3_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_3_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_3_io_in_stage = local_pes_20_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_4_clock = clock;
  assign local_pes_20_4_reset = reset;
  assign local_pes_20_4_io_in_q = local_pes_20_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_4_io_in_sum = local_pes_20_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_4_io_in_sum_exp = local_pes_20_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_4_io_in_kv = local_pes_19_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_4_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_4_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_4_io_in_stage = local_pes_20_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_5_clock = clock;
  assign local_pes_20_5_reset = reset;
  assign local_pes_20_5_io_in_q = local_pes_20_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_5_io_in_sum = local_pes_20_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_5_io_in_sum_exp = local_pes_20_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_5_io_in_kv = local_pes_19_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_5_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_5_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_5_io_in_stage = local_pes_20_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_6_clock = clock;
  assign local_pes_20_6_reset = reset;
  assign local_pes_20_6_io_in_q = local_pes_20_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_6_io_in_sum = local_pes_20_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_6_io_in_sum_exp = local_pes_20_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_6_io_in_kv = local_pes_19_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_6_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_6_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_6_io_in_stage = local_pes_20_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_7_clock = clock;
  assign local_pes_20_7_reset = reset;
  assign local_pes_20_7_io_in_q = local_pes_20_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_7_io_in_sum = local_pes_20_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_7_io_in_sum_exp = local_pes_20_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_7_io_in_kv = local_pes_19_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_7_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_7_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_7_io_in_stage = local_pes_20_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_8_clock = clock;
  assign local_pes_20_8_reset = reset;
  assign local_pes_20_8_io_in_q = local_pes_20_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_8_io_in_sum = local_pes_20_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_8_io_in_sum_exp = local_pes_20_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_8_io_in_kv = local_pes_19_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_8_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_8_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_8_io_in_stage = local_pes_20_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_9_clock = clock;
  assign local_pes_20_9_reset = reset;
  assign local_pes_20_9_io_in_q = local_pes_20_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_9_io_in_sum = local_pes_20_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_9_io_in_sum_exp = local_pes_20_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_9_io_in_kv = local_pes_19_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_9_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_9_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_9_io_in_stage = local_pes_20_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_10_clock = clock;
  assign local_pes_20_10_reset = reset;
  assign local_pes_20_10_io_in_q = local_pes_20_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_10_io_in_sum = local_pes_20_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_10_io_in_sum_exp = local_pes_20_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_10_io_in_kv = local_pes_19_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_10_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_10_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_10_io_in_stage = local_pes_20_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_11_clock = clock;
  assign local_pes_20_11_reset = reset;
  assign local_pes_20_11_io_in_q = local_pes_20_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_11_io_in_sum = local_pes_20_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_11_io_in_sum_exp = local_pes_20_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_11_io_in_kv = local_pes_19_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_11_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_11_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_11_io_in_stage = local_pes_20_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_12_clock = clock;
  assign local_pes_20_12_reset = reset;
  assign local_pes_20_12_io_in_q = local_pes_20_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_12_io_in_sum = local_pes_20_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_12_io_in_sum_exp = local_pes_20_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_12_io_in_kv = local_pes_19_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_12_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_12_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_12_io_in_stage = local_pes_20_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_13_clock = clock;
  assign local_pes_20_13_reset = reset;
  assign local_pes_20_13_io_in_q = local_pes_20_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_13_io_in_sum = local_pes_20_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_13_io_in_sum_exp = local_pes_20_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_13_io_in_kv = local_pes_19_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_13_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_13_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_13_io_in_stage = local_pes_20_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_14_clock = clock;
  assign local_pes_20_14_reset = reset;
  assign local_pes_20_14_io_in_q = local_pes_20_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_14_io_in_sum = local_pes_20_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_14_io_in_sum_exp = local_pes_20_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_14_io_in_kv = local_pes_19_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_14_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_14_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_14_io_in_stage = local_pes_20_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_15_clock = clock;
  assign local_pes_20_15_reset = reset;
  assign local_pes_20_15_io_in_q = local_pes_20_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_15_io_in_sum = local_pes_20_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_15_io_in_sum_exp = local_pes_20_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_15_io_in_kv = local_pes_19_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_15_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_15_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_15_io_in_stage = local_pes_20_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_16_clock = clock;
  assign local_pes_20_16_reset = reset;
  assign local_pes_20_16_io_in_q = local_pes_20_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_16_io_in_sum = local_pes_20_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_16_io_in_sum_exp = local_pes_20_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_16_io_in_kv = local_pes_19_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_16_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_16_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_16_io_in_stage = local_pes_20_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_17_clock = clock;
  assign local_pes_20_17_reset = reset;
  assign local_pes_20_17_io_in_q = local_pes_20_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_17_io_in_sum = local_pes_20_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_17_io_in_sum_exp = local_pes_20_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_17_io_in_kv = local_pes_19_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_17_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_17_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_17_io_in_stage = local_pes_20_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_18_clock = clock;
  assign local_pes_20_18_reset = reset;
  assign local_pes_20_18_io_in_q = local_pes_20_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_18_io_in_sum = local_pes_20_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_18_io_in_sum_exp = local_pes_20_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_18_io_in_kv = local_pes_19_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_18_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_18_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_18_io_in_stage = local_pes_20_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_19_clock = clock;
  assign local_pes_20_19_reset = reset;
  assign local_pes_20_19_io_in_q = local_pes_20_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_19_io_in_sum = local_pes_20_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_19_io_in_sum_exp = local_pes_20_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_19_io_in_kv = local_pes_19_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_19_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_19_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_19_io_in_stage = local_pes_20_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_20_clock = clock;
  assign local_pes_20_20_reset = reset;
  assign local_pes_20_20_io_in_q = local_pes_20_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_20_io_in_sum = local_pes_20_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_20_io_in_sum_exp = local_pes_20_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_20_io_in_kv = local_pes_19_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_20_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_20_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_20_io_in_stage = local_pes_20_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_21_clock = clock;
  assign local_pes_20_21_reset = reset;
  assign local_pes_20_21_io_in_q = local_pes_20_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_21_io_in_sum = local_pes_20_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_21_io_in_sum_exp = local_pes_20_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_21_io_in_kv = local_pes_19_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_21_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_21_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_21_io_in_stage = local_pes_20_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_22_clock = clock;
  assign local_pes_20_22_reset = reset;
  assign local_pes_20_22_io_in_q = local_pes_20_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_22_io_in_sum = local_pes_20_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_22_io_in_sum_exp = local_pes_20_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_22_io_in_kv = local_pes_19_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_22_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_22_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_22_io_in_stage = local_pes_20_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_23_clock = clock;
  assign local_pes_20_23_reset = reset;
  assign local_pes_20_23_io_in_q = local_pes_20_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_23_io_in_sum = local_pes_20_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_23_io_in_sum_exp = local_pes_20_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_23_io_in_kv = local_pes_19_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_23_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_23_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_23_io_in_stage = local_pes_20_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_24_clock = clock;
  assign local_pes_20_24_reset = reset;
  assign local_pes_20_24_io_in_q = local_pes_20_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_24_io_in_sum = local_pes_20_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_24_io_in_sum_exp = local_pes_20_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_24_io_in_kv = local_pes_19_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_24_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_24_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_24_io_in_stage = local_pes_20_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_25_clock = clock;
  assign local_pes_20_25_reset = reset;
  assign local_pes_20_25_io_in_q = local_pes_20_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_25_io_in_sum = local_pes_20_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_25_io_in_sum_exp = local_pes_20_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_25_io_in_kv = local_pes_19_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_25_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_25_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_25_io_in_stage = local_pes_20_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_26_clock = clock;
  assign local_pes_20_26_reset = reset;
  assign local_pes_20_26_io_in_q = local_pes_20_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_26_io_in_sum = local_pes_20_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_26_io_in_sum_exp = local_pes_20_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_26_io_in_kv = local_pes_19_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_26_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_26_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_26_io_in_stage = local_pes_20_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_27_clock = clock;
  assign local_pes_20_27_reset = reset;
  assign local_pes_20_27_io_in_q = local_pes_20_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_27_io_in_sum = local_pes_20_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_27_io_in_sum_exp = local_pes_20_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_27_io_in_kv = local_pes_19_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_27_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_27_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_27_io_in_stage = local_pes_20_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_28_clock = clock;
  assign local_pes_20_28_reset = reset;
  assign local_pes_20_28_io_in_q = local_pes_20_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_28_io_in_sum = local_pes_20_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_28_io_in_sum_exp = local_pes_20_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_28_io_in_kv = local_pes_19_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_28_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_28_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_28_io_in_stage = local_pes_20_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_29_clock = clock;
  assign local_pes_20_29_reset = reset;
  assign local_pes_20_29_io_in_q = local_pes_20_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_29_io_in_sum = local_pes_20_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_29_io_in_sum_exp = local_pes_20_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_29_io_in_kv = local_pes_19_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_29_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_29_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_29_io_in_stage = local_pes_20_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_30_clock = clock;
  assign local_pes_20_30_reset = reset;
  assign local_pes_20_30_io_in_q = local_pes_20_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_30_io_in_sum = local_pes_20_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_30_io_in_sum_exp = local_pes_20_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_30_io_in_kv = local_pes_19_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_30_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_30_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_30_io_in_stage = local_pes_20_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_20_31_clock = clock;
  assign local_pes_20_31_reset = reset;
  assign local_pes_20_31_io_in_q = local_pes_20_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_20_31_io_in_sum = local_pes_20_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_20_31_io_in_sum_exp = local_pes_20_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_20_31_io_in_kv = local_pes_19_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_20_31_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_20_31_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_20_31_io_in_stage = local_pes_20_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_0_clock = clock;
  assign local_pes_21_0_reset = reset;
  assign local_pes_21_0_io_in_q = io_q_ports_21; // @[PEArray.scala 51:37]
  assign local_pes_21_0_io_in_kv = io_kv_ports_52; // @[PEArray.scala 40:34]
  assign local_pes_21_0_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_0_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_0_io_in_stage = io_stage_ports_21; // @[PEArray.scala 52:41]
  assign local_pes_21_1_clock = clock;
  assign local_pes_21_1_reset = reset;
  assign local_pes_21_1_io_in_q = local_pes_21_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_1_io_in_sum = local_pes_21_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_21_1_io_in_kv = local_pes_20_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_1_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_1_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_1_io_in_stage = local_pes_21_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_2_clock = clock;
  assign local_pes_21_2_reset = reset;
  assign local_pes_21_2_io_in_q = local_pes_21_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_2_io_in_sum = local_pes_21_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_2_io_in_sum_exp = local_pes_21_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_2_io_in_kv = local_pes_20_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_2_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_2_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_2_io_in_stage = local_pes_21_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_3_clock = clock;
  assign local_pes_21_3_reset = reset;
  assign local_pes_21_3_io_in_q = local_pes_21_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_3_io_in_sum = local_pes_21_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_3_io_in_sum_exp = local_pes_21_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_3_io_in_kv = local_pes_20_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_3_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_3_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_3_io_in_stage = local_pes_21_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_4_clock = clock;
  assign local_pes_21_4_reset = reset;
  assign local_pes_21_4_io_in_q = local_pes_21_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_4_io_in_sum = local_pes_21_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_4_io_in_sum_exp = local_pes_21_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_4_io_in_kv = local_pes_20_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_4_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_4_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_4_io_in_stage = local_pes_21_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_5_clock = clock;
  assign local_pes_21_5_reset = reset;
  assign local_pes_21_5_io_in_q = local_pes_21_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_5_io_in_sum = local_pes_21_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_5_io_in_sum_exp = local_pes_21_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_5_io_in_kv = local_pes_20_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_5_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_5_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_5_io_in_stage = local_pes_21_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_6_clock = clock;
  assign local_pes_21_6_reset = reset;
  assign local_pes_21_6_io_in_q = local_pes_21_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_6_io_in_sum = local_pes_21_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_6_io_in_sum_exp = local_pes_21_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_6_io_in_kv = local_pes_20_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_6_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_6_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_6_io_in_stage = local_pes_21_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_7_clock = clock;
  assign local_pes_21_7_reset = reset;
  assign local_pes_21_7_io_in_q = local_pes_21_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_7_io_in_sum = local_pes_21_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_7_io_in_sum_exp = local_pes_21_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_7_io_in_kv = local_pes_20_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_7_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_7_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_7_io_in_stage = local_pes_21_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_8_clock = clock;
  assign local_pes_21_8_reset = reset;
  assign local_pes_21_8_io_in_q = local_pes_21_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_8_io_in_sum = local_pes_21_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_8_io_in_sum_exp = local_pes_21_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_8_io_in_kv = local_pes_20_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_8_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_8_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_8_io_in_stage = local_pes_21_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_9_clock = clock;
  assign local_pes_21_9_reset = reset;
  assign local_pes_21_9_io_in_q = local_pes_21_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_9_io_in_sum = local_pes_21_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_9_io_in_sum_exp = local_pes_21_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_9_io_in_kv = local_pes_20_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_9_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_9_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_9_io_in_stage = local_pes_21_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_10_clock = clock;
  assign local_pes_21_10_reset = reset;
  assign local_pes_21_10_io_in_q = local_pes_21_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_10_io_in_sum = local_pes_21_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_10_io_in_sum_exp = local_pes_21_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_10_io_in_kv = local_pes_20_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_10_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_10_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_10_io_in_stage = local_pes_21_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_11_clock = clock;
  assign local_pes_21_11_reset = reset;
  assign local_pes_21_11_io_in_q = local_pes_21_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_11_io_in_sum = local_pes_21_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_11_io_in_sum_exp = local_pes_21_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_11_io_in_kv = local_pes_20_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_11_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_11_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_11_io_in_stage = local_pes_21_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_12_clock = clock;
  assign local_pes_21_12_reset = reset;
  assign local_pes_21_12_io_in_q = local_pes_21_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_12_io_in_sum = local_pes_21_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_12_io_in_sum_exp = local_pes_21_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_12_io_in_kv = local_pes_20_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_12_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_12_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_12_io_in_stage = local_pes_21_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_13_clock = clock;
  assign local_pes_21_13_reset = reset;
  assign local_pes_21_13_io_in_q = local_pes_21_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_13_io_in_sum = local_pes_21_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_13_io_in_sum_exp = local_pes_21_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_13_io_in_kv = local_pes_20_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_13_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_13_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_13_io_in_stage = local_pes_21_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_14_clock = clock;
  assign local_pes_21_14_reset = reset;
  assign local_pes_21_14_io_in_q = local_pes_21_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_14_io_in_sum = local_pes_21_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_14_io_in_sum_exp = local_pes_21_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_14_io_in_kv = local_pes_20_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_14_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_14_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_14_io_in_stage = local_pes_21_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_15_clock = clock;
  assign local_pes_21_15_reset = reset;
  assign local_pes_21_15_io_in_q = local_pes_21_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_15_io_in_sum = local_pes_21_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_15_io_in_sum_exp = local_pes_21_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_15_io_in_kv = local_pes_20_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_15_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_15_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_15_io_in_stage = local_pes_21_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_16_clock = clock;
  assign local_pes_21_16_reset = reset;
  assign local_pes_21_16_io_in_q = local_pes_21_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_16_io_in_sum = local_pes_21_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_16_io_in_sum_exp = local_pes_21_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_16_io_in_kv = local_pes_20_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_16_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_16_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_16_io_in_stage = local_pes_21_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_17_clock = clock;
  assign local_pes_21_17_reset = reset;
  assign local_pes_21_17_io_in_q = local_pes_21_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_17_io_in_sum = local_pes_21_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_17_io_in_sum_exp = local_pes_21_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_17_io_in_kv = local_pes_20_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_17_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_17_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_17_io_in_stage = local_pes_21_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_18_clock = clock;
  assign local_pes_21_18_reset = reset;
  assign local_pes_21_18_io_in_q = local_pes_21_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_18_io_in_sum = local_pes_21_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_18_io_in_sum_exp = local_pes_21_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_18_io_in_kv = local_pes_20_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_18_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_18_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_18_io_in_stage = local_pes_21_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_19_clock = clock;
  assign local_pes_21_19_reset = reset;
  assign local_pes_21_19_io_in_q = local_pes_21_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_19_io_in_sum = local_pes_21_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_19_io_in_sum_exp = local_pes_21_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_19_io_in_kv = local_pes_20_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_19_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_19_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_19_io_in_stage = local_pes_21_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_20_clock = clock;
  assign local_pes_21_20_reset = reset;
  assign local_pes_21_20_io_in_q = local_pes_21_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_20_io_in_sum = local_pes_21_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_20_io_in_sum_exp = local_pes_21_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_20_io_in_kv = local_pes_20_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_20_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_20_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_20_io_in_stage = local_pes_21_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_21_clock = clock;
  assign local_pes_21_21_reset = reset;
  assign local_pes_21_21_io_in_q = local_pes_21_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_21_io_in_sum = local_pes_21_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_21_io_in_sum_exp = local_pes_21_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_21_io_in_kv = local_pes_20_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_21_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_21_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_21_io_in_stage = local_pes_21_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_22_clock = clock;
  assign local_pes_21_22_reset = reset;
  assign local_pes_21_22_io_in_q = local_pes_21_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_22_io_in_sum = local_pes_21_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_22_io_in_sum_exp = local_pes_21_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_22_io_in_kv = local_pes_20_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_22_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_22_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_22_io_in_stage = local_pes_21_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_23_clock = clock;
  assign local_pes_21_23_reset = reset;
  assign local_pes_21_23_io_in_q = local_pes_21_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_23_io_in_sum = local_pes_21_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_23_io_in_sum_exp = local_pes_21_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_23_io_in_kv = local_pes_20_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_23_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_23_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_23_io_in_stage = local_pes_21_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_24_clock = clock;
  assign local_pes_21_24_reset = reset;
  assign local_pes_21_24_io_in_q = local_pes_21_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_24_io_in_sum = local_pes_21_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_24_io_in_sum_exp = local_pes_21_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_24_io_in_kv = local_pes_20_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_24_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_24_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_24_io_in_stage = local_pes_21_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_25_clock = clock;
  assign local_pes_21_25_reset = reset;
  assign local_pes_21_25_io_in_q = local_pes_21_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_25_io_in_sum = local_pes_21_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_25_io_in_sum_exp = local_pes_21_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_25_io_in_kv = local_pes_20_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_25_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_25_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_25_io_in_stage = local_pes_21_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_26_clock = clock;
  assign local_pes_21_26_reset = reset;
  assign local_pes_21_26_io_in_q = local_pes_21_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_26_io_in_sum = local_pes_21_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_26_io_in_sum_exp = local_pes_21_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_26_io_in_kv = local_pes_20_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_26_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_26_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_26_io_in_stage = local_pes_21_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_27_clock = clock;
  assign local_pes_21_27_reset = reset;
  assign local_pes_21_27_io_in_q = local_pes_21_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_27_io_in_sum = local_pes_21_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_27_io_in_sum_exp = local_pes_21_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_27_io_in_kv = local_pes_20_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_27_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_27_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_27_io_in_stage = local_pes_21_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_28_clock = clock;
  assign local_pes_21_28_reset = reset;
  assign local_pes_21_28_io_in_q = local_pes_21_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_28_io_in_sum = local_pes_21_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_28_io_in_sum_exp = local_pes_21_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_28_io_in_kv = local_pes_20_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_28_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_28_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_28_io_in_stage = local_pes_21_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_29_clock = clock;
  assign local_pes_21_29_reset = reset;
  assign local_pes_21_29_io_in_q = local_pes_21_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_29_io_in_sum = local_pes_21_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_29_io_in_sum_exp = local_pes_21_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_29_io_in_kv = local_pes_20_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_29_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_29_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_29_io_in_stage = local_pes_21_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_30_clock = clock;
  assign local_pes_21_30_reset = reset;
  assign local_pes_21_30_io_in_q = local_pes_21_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_30_io_in_sum = local_pes_21_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_30_io_in_sum_exp = local_pes_21_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_30_io_in_kv = local_pes_20_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_30_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_30_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_30_io_in_stage = local_pes_21_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_21_31_clock = clock;
  assign local_pes_21_31_reset = reset;
  assign local_pes_21_31_io_in_q = local_pes_21_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_21_31_io_in_sum = local_pes_21_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_21_31_io_in_sum_exp = local_pes_21_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_21_31_io_in_kv = local_pes_20_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_21_31_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_21_31_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_21_31_io_in_stage = local_pes_21_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_0_clock = clock;
  assign local_pes_22_0_reset = reset;
  assign local_pes_22_0_io_in_q = io_q_ports_22; // @[PEArray.scala 51:37]
  assign local_pes_22_0_io_in_kv = io_kv_ports_53; // @[PEArray.scala 40:34]
  assign local_pes_22_0_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_0_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_0_io_in_stage = io_stage_ports_22; // @[PEArray.scala 52:41]
  assign local_pes_22_1_clock = clock;
  assign local_pes_22_1_reset = reset;
  assign local_pes_22_1_io_in_q = local_pes_22_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_1_io_in_sum = local_pes_22_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_22_1_io_in_kv = local_pes_21_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_1_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_1_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_1_io_in_stage = local_pes_22_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_2_clock = clock;
  assign local_pes_22_2_reset = reset;
  assign local_pes_22_2_io_in_q = local_pes_22_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_2_io_in_sum = local_pes_22_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_2_io_in_sum_exp = local_pes_22_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_2_io_in_kv = local_pes_21_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_2_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_2_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_2_io_in_stage = local_pes_22_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_3_clock = clock;
  assign local_pes_22_3_reset = reset;
  assign local_pes_22_3_io_in_q = local_pes_22_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_3_io_in_sum = local_pes_22_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_3_io_in_sum_exp = local_pes_22_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_3_io_in_kv = local_pes_21_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_3_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_3_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_3_io_in_stage = local_pes_22_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_4_clock = clock;
  assign local_pes_22_4_reset = reset;
  assign local_pes_22_4_io_in_q = local_pes_22_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_4_io_in_sum = local_pes_22_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_4_io_in_sum_exp = local_pes_22_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_4_io_in_kv = local_pes_21_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_4_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_4_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_4_io_in_stage = local_pes_22_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_5_clock = clock;
  assign local_pes_22_5_reset = reset;
  assign local_pes_22_5_io_in_q = local_pes_22_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_5_io_in_sum = local_pes_22_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_5_io_in_sum_exp = local_pes_22_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_5_io_in_kv = local_pes_21_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_5_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_5_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_5_io_in_stage = local_pes_22_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_6_clock = clock;
  assign local_pes_22_6_reset = reset;
  assign local_pes_22_6_io_in_q = local_pes_22_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_6_io_in_sum = local_pes_22_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_6_io_in_sum_exp = local_pes_22_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_6_io_in_kv = local_pes_21_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_6_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_6_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_6_io_in_stage = local_pes_22_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_7_clock = clock;
  assign local_pes_22_7_reset = reset;
  assign local_pes_22_7_io_in_q = local_pes_22_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_7_io_in_sum = local_pes_22_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_7_io_in_sum_exp = local_pes_22_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_7_io_in_kv = local_pes_21_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_7_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_7_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_7_io_in_stage = local_pes_22_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_8_clock = clock;
  assign local_pes_22_8_reset = reset;
  assign local_pes_22_8_io_in_q = local_pes_22_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_8_io_in_sum = local_pes_22_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_8_io_in_sum_exp = local_pes_22_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_8_io_in_kv = local_pes_21_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_8_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_8_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_8_io_in_stage = local_pes_22_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_9_clock = clock;
  assign local_pes_22_9_reset = reset;
  assign local_pes_22_9_io_in_q = local_pes_22_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_9_io_in_sum = local_pes_22_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_9_io_in_sum_exp = local_pes_22_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_9_io_in_kv = local_pes_21_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_9_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_9_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_9_io_in_stage = local_pes_22_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_10_clock = clock;
  assign local_pes_22_10_reset = reset;
  assign local_pes_22_10_io_in_q = local_pes_22_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_10_io_in_sum = local_pes_22_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_10_io_in_sum_exp = local_pes_22_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_10_io_in_kv = local_pes_21_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_10_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_10_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_10_io_in_stage = local_pes_22_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_11_clock = clock;
  assign local_pes_22_11_reset = reset;
  assign local_pes_22_11_io_in_q = local_pes_22_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_11_io_in_sum = local_pes_22_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_11_io_in_sum_exp = local_pes_22_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_11_io_in_kv = local_pes_21_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_11_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_11_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_11_io_in_stage = local_pes_22_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_12_clock = clock;
  assign local_pes_22_12_reset = reset;
  assign local_pes_22_12_io_in_q = local_pes_22_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_12_io_in_sum = local_pes_22_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_12_io_in_sum_exp = local_pes_22_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_12_io_in_kv = local_pes_21_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_12_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_12_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_12_io_in_stage = local_pes_22_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_13_clock = clock;
  assign local_pes_22_13_reset = reset;
  assign local_pes_22_13_io_in_q = local_pes_22_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_13_io_in_sum = local_pes_22_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_13_io_in_sum_exp = local_pes_22_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_13_io_in_kv = local_pes_21_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_13_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_13_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_13_io_in_stage = local_pes_22_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_14_clock = clock;
  assign local_pes_22_14_reset = reset;
  assign local_pes_22_14_io_in_q = local_pes_22_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_14_io_in_sum = local_pes_22_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_14_io_in_sum_exp = local_pes_22_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_14_io_in_kv = local_pes_21_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_14_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_14_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_14_io_in_stage = local_pes_22_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_15_clock = clock;
  assign local_pes_22_15_reset = reset;
  assign local_pes_22_15_io_in_q = local_pes_22_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_15_io_in_sum = local_pes_22_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_15_io_in_sum_exp = local_pes_22_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_15_io_in_kv = local_pes_21_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_15_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_15_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_15_io_in_stage = local_pes_22_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_16_clock = clock;
  assign local_pes_22_16_reset = reset;
  assign local_pes_22_16_io_in_q = local_pes_22_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_16_io_in_sum = local_pes_22_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_16_io_in_sum_exp = local_pes_22_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_16_io_in_kv = local_pes_21_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_16_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_16_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_16_io_in_stage = local_pes_22_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_17_clock = clock;
  assign local_pes_22_17_reset = reset;
  assign local_pes_22_17_io_in_q = local_pes_22_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_17_io_in_sum = local_pes_22_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_17_io_in_sum_exp = local_pes_22_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_17_io_in_kv = local_pes_21_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_17_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_17_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_17_io_in_stage = local_pes_22_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_18_clock = clock;
  assign local_pes_22_18_reset = reset;
  assign local_pes_22_18_io_in_q = local_pes_22_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_18_io_in_sum = local_pes_22_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_18_io_in_sum_exp = local_pes_22_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_18_io_in_kv = local_pes_21_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_18_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_18_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_18_io_in_stage = local_pes_22_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_19_clock = clock;
  assign local_pes_22_19_reset = reset;
  assign local_pes_22_19_io_in_q = local_pes_22_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_19_io_in_sum = local_pes_22_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_19_io_in_sum_exp = local_pes_22_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_19_io_in_kv = local_pes_21_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_19_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_19_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_19_io_in_stage = local_pes_22_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_20_clock = clock;
  assign local_pes_22_20_reset = reset;
  assign local_pes_22_20_io_in_q = local_pes_22_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_20_io_in_sum = local_pes_22_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_20_io_in_sum_exp = local_pes_22_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_20_io_in_kv = local_pes_21_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_20_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_20_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_20_io_in_stage = local_pes_22_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_21_clock = clock;
  assign local_pes_22_21_reset = reset;
  assign local_pes_22_21_io_in_q = local_pes_22_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_21_io_in_sum = local_pes_22_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_21_io_in_sum_exp = local_pes_22_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_21_io_in_kv = local_pes_21_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_21_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_21_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_21_io_in_stage = local_pes_22_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_22_clock = clock;
  assign local_pes_22_22_reset = reset;
  assign local_pes_22_22_io_in_q = local_pes_22_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_22_io_in_sum = local_pes_22_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_22_io_in_sum_exp = local_pes_22_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_22_io_in_kv = local_pes_21_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_22_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_22_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_22_io_in_stage = local_pes_22_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_23_clock = clock;
  assign local_pes_22_23_reset = reset;
  assign local_pes_22_23_io_in_q = local_pes_22_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_23_io_in_sum = local_pes_22_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_23_io_in_sum_exp = local_pes_22_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_23_io_in_kv = local_pes_21_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_23_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_23_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_23_io_in_stage = local_pes_22_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_24_clock = clock;
  assign local_pes_22_24_reset = reset;
  assign local_pes_22_24_io_in_q = local_pes_22_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_24_io_in_sum = local_pes_22_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_24_io_in_sum_exp = local_pes_22_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_24_io_in_kv = local_pes_21_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_24_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_24_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_24_io_in_stage = local_pes_22_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_25_clock = clock;
  assign local_pes_22_25_reset = reset;
  assign local_pes_22_25_io_in_q = local_pes_22_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_25_io_in_sum = local_pes_22_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_25_io_in_sum_exp = local_pes_22_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_25_io_in_kv = local_pes_21_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_25_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_25_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_25_io_in_stage = local_pes_22_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_26_clock = clock;
  assign local_pes_22_26_reset = reset;
  assign local_pes_22_26_io_in_q = local_pes_22_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_26_io_in_sum = local_pes_22_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_26_io_in_sum_exp = local_pes_22_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_26_io_in_kv = local_pes_21_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_26_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_26_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_26_io_in_stage = local_pes_22_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_27_clock = clock;
  assign local_pes_22_27_reset = reset;
  assign local_pes_22_27_io_in_q = local_pes_22_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_27_io_in_sum = local_pes_22_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_27_io_in_sum_exp = local_pes_22_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_27_io_in_kv = local_pes_21_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_27_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_27_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_27_io_in_stage = local_pes_22_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_28_clock = clock;
  assign local_pes_22_28_reset = reset;
  assign local_pes_22_28_io_in_q = local_pes_22_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_28_io_in_sum = local_pes_22_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_28_io_in_sum_exp = local_pes_22_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_28_io_in_kv = local_pes_21_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_28_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_28_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_28_io_in_stage = local_pes_22_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_29_clock = clock;
  assign local_pes_22_29_reset = reset;
  assign local_pes_22_29_io_in_q = local_pes_22_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_29_io_in_sum = local_pes_22_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_29_io_in_sum_exp = local_pes_22_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_29_io_in_kv = local_pes_21_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_29_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_29_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_29_io_in_stage = local_pes_22_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_30_clock = clock;
  assign local_pes_22_30_reset = reset;
  assign local_pes_22_30_io_in_q = local_pes_22_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_30_io_in_sum = local_pes_22_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_30_io_in_sum_exp = local_pes_22_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_30_io_in_kv = local_pes_21_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_30_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_30_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_30_io_in_stage = local_pes_22_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_22_31_clock = clock;
  assign local_pes_22_31_reset = reset;
  assign local_pes_22_31_io_in_q = local_pes_22_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_22_31_io_in_sum = local_pes_22_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_22_31_io_in_sum_exp = local_pes_22_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_22_31_io_in_kv = local_pes_21_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_22_31_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_22_31_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_22_31_io_in_stage = local_pes_22_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_0_clock = clock;
  assign local_pes_23_0_reset = reset;
  assign local_pes_23_0_io_in_q = io_q_ports_23; // @[PEArray.scala 51:37]
  assign local_pes_23_0_io_in_kv = io_kv_ports_54; // @[PEArray.scala 40:34]
  assign local_pes_23_0_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_0_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_0_io_in_stage = io_stage_ports_23; // @[PEArray.scala 52:41]
  assign local_pes_23_1_clock = clock;
  assign local_pes_23_1_reset = reset;
  assign local_pes_23_1_io_in_q = local_pes_23_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_1_io_in_sum = local_pes_23_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_23_1_io_in_kv = local_pes_22_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_1_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_1_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_1_io_in_stage = local_pes_23_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_2_clock = clock;
  assign local_pes_23_2_reset = reset;
  assign local_pes_23_2_io_in_q = local_pes_23_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_2_io_in_sum = local_pes_23_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_2_io_in_sum_exp = local_pes_23_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_2_io_in_kv = local_pes_22_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_2_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_2_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_2_io_in_stage = local_pes_23_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_3_clock = clock;
  assign local_pes_23_3_reset = reset;
  assign local_pes_23_3_io_in_q = local_pes_23_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_3_io_in_sum = local_pes_23_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_3_io_in_sum_exp = local_pes_23_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_3_io_in_kv = local_pes_22_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_3_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_3_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_3_io_in_stage = local_pes_23_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_4_clock = clock;
  assign local_pes_23_4_reset = reset;
  assign local_pes_23_4_io_in_q = local_pes_23_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_4_io_in_sum = local_pes_23_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_4_io_in_sum_exp = local_pes_23_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_4_io_in_kv = local_pes_22_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_4_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_4_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_4_io_in_stage = local_pes_23_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_5_clock = clock;
  assign local_pes_23_5_reset = reset;
  assign local_pes_23_5_io_in_q = local_pes_23_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_5_io_in_sum = local_pes_23_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_5_io_in_sum_exp = local_pes_23_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_5_io_in_kv = local_pes_22_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_5_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_5_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_5_io_in_stage = local_pes_23_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_6_clock = clock;
  assign local_pes_23_6_reset = reset;
  assign local_pes_23_6_io_in_q = local_pes_23_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_6_io_in_sum = local_pes_23_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_6_io_in_sum_exp = local_pes_23_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_6_io_in_kv = local_pes_22_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_6_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_6_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_6_io_in_stage = local_pes_23_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_7_clock = clock;
  assign local_pes_23_7_reset = reset;
  assign local_pes_23_7_io_in_q = local_pes_23_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_7_io_in_sum = local_pes_23_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_7_io_in_sum_exp = local_pes_23_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_7_io_in_kv = local_pes_22_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_7_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_7_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_7_io_in_stage = local_pes_23_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_8_clock = clock;
  assign local_pes_23_8_reset = reset;
  assign local_pes_23_8_io_in_q = local_pes_23_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_8_io_in_sum = local_pes_23_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_8_io_in_sum_exp = local_pes_23_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_8_io_in_kv = local_pes_22_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_8_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_8_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_8_io_in_stage = local_pes_23_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_9_clock = clock;
  assign local_pes_23_9_reset = reset;
  assign local_pes_23_9_io_in_q = local_pes_23_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_9_io_in_sum = local_pes_23_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_9_io_in_sum_exp = local_pes_23_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_9_io_in_kv = local_pes_22_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_9_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_9_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_9_io_in_stage = local_pes_23_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_10_clock = clock;
  assign local_pes_23_10_reset = reset;
  assign local_pes_23_10_io_in_q = local_pes_23_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_10_io_in_sum = local_pes_23_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_10_io_in_sum_exp = local_pes_23_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_10_io_in_kv = local_pes_22_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_10_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_10_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_10_io_in_stage = local_pes_23_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_11_clock = clock;
  assign local_pes_23_11_reset = reset;
  assign local_pes_23_11_io_in_q = local_pes_23_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_11_io_in_sum = local_pes_23_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_11_io_in_sum_exp = local_pes_23_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_11_io_in_kv = local_pes_22_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_11_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_11_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_11_io_in_stage = local_pes_23_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_12_clock = clock;
  assign local_pes_23_12_reset = reset;
  assign local_pes_23_12_io_in_q = local_pes_23_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_12_io_in_sum = local_pes_23_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_12_io_in_sum_exp = local_pes_23_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_12_io_in_kv = local_pes_22_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_12_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_12_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_12_io_in_stage = local_pes_23_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_13_clock = clock;
  assign local_pes_23_13_reset = reset;
  assign local_pes_23_13_io_in_q = local_pes_23_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_13_io_in_sum = local_pes_23_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_13_io_in_sum_exp = local_pes_23_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_13_io_in_kv = local_pes_22_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_13_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_13_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_13_io_in_stage = local_pes_23_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_14_clock = clock;
  assign local_pes_23_14_reset = reset;
  assign local_pes_23_14_io_in_q = local_pes_23_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_14_io_in_sum = local_pes_23_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_14_io_in_sum_exp = local_pes_23_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_14_io_in_kv = local_pes_22_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_14_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_14_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_14_io_in_stage = local_pes_23_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_15_clock = clock;
  assign local_pes_23_15_reset = reset;
  assign local_pes_23_15_io_in_q = local_pes_23_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_15_io_in_sum = local_pes_23_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_15_io_in_sum_exp = local_pes_23_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_15_io_in_kv = local_pes_22_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_15_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_15_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_15_io_in_stage = local_pes_23_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_16_clock = clock;
  assign local_pes_23_16_reset = reset;
  assign local_pes_23_16_io_in_q = local_pes_23_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_16_io_in_sum = local_pes_23_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_16_io_in_sum_exp = local_pes_23_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_16_io_in_kv = local_pes_22_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_16_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_16_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_16_io_in_stage = local_pes_23_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_17_clock = clock;
  assign local_pes_23_17_reset = reset;
  assign local_pes_23_17_io_in_q = local_pes_23_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_17_io_in_sum = local_pes_23_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_17_io_in_sum_exp = local_pes_23_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_17_io_in_kv = local_pes_22_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_17_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_17_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_17_io_in_stage = local_pes_23_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_18_clock = clock;
  assign local_pes_23_18_reset = reset;
  assign local_pes_23_18_io_in_q = local_pes_23_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_18_io_in_sum = local_pes_23_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_18_io_in_sum_exp = local_pes_23_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_18_io_in_kv = local_pes_22_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_18_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_18_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_18_io_in_stage = local_pes_23_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_19_clock = clock;
  assign local_pes_23_19_reset = reset;
  assign local_pes_23_19_io_in_q = local_pes_23_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_19_io_in_sum = local_pes_23_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_19_io_in_sum_exp = local_pes_23_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_19_io_in_kv = local_pes_22_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_19_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_19_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_19_io_in_stage = local_pes_23_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_20_clock = clock;
  assign local_pes_23_20_reset = reset;
  assign local_pes_23_20_io_in_q = local_pes_23_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_20_io_in_sum = local_pes_23_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_20_io_in_sum_exp = local_pes_23_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_20_io_in_kv = local_pes_22_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_20_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_20_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_20_io_in_stage = local_pes_23_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_21_clock = clock;
  assign local_pes_23_21_reset = reset;
  assign local_pes_23_21_io_in_q = local_pes_23_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_21_io_in_sum = local_pes_23_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_21_io_in_sum_exp = local_pes_23_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_21_io_in_kv = local_pes_22_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_21_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_21_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_21_io_in_stage = local_pes_23_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_22_clock = clock;
  assign local_pes_23_22_reset = reset;
  assign local_pes_23_22_io_in_q = local_pes_23_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_22_io_in_sum = local_pes_23_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_22_io_in_sum_exp = local_pes_23_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_22_io_in_kv = local_pes_22_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_22_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_22_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_22_io_in_stage = local_pes_23_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_23_clock = clock;
  assign local_pes_23_23_reset = reset;
  assign local_pes_23_23_io_in_q = local_pes_23_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_23_io_in_sum = local_pes_23_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_23_io_in_sum_exp = local_pes_23_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_23_io_in_kv = local_pes_22_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_23_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_23_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_23_io_in_stage = local_pes_23_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_24_clock = clock;
  assign local_pes_23_24_reset = reset;
  assign local_pes_23_24_io_in_q = local_pes_23_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_24_io_in_sum = local_pes_23_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_24_io_in_sum_exp = local_pes_23_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_24_io_in_kv = local_pes_22_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_24_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_24_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_24_io_in_stage = local_pes_23_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_25_clock = clock;
  assign local_pes_23_25_reset = reset;
  assign local_pes_23_25_io_in_q = local_pes_23_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_25_io_in_sum = local_pes_23_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_25_io_in_sum_exp = local_pes_23_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_25_io_in_kv = local_pes_22_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_25_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_25_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_25_io_in_stage = local_pes_23_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_26_clock = clock;
  assign local_pes_23_26_reset = reset;
  assign local_pes_23_26_io_in_q = local_pes_23_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_26_io_in_sum = local_pes_23_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_26_io_in_sum_exp = local_pes_23_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_26_io_in_kv = local_pes_22_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_26_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_26_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_26_io_in_stage = local_pes_23_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_27_clock = clock;
  assign local_pes_23_27_reset = reset;
  assign local_pes_23_27_io_in_q = local_pes_23_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_27_io_in_sum = local_pes_23_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_27_io_in_sum_exp = local_pes_23_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_27_io_in_kv = local_pes_22_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_27_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_27_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_27_io_in_stage = local_pes_23_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_28_clock = clock;
  assign local_pes_23_28_reset = reset;
  assign local_pes_23_28_io_in_q = local_pes_23_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_28_io_in_sum = local_pes_23_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_28_io_in_sum_exp = local_pes_23_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_28_io_in_kv = local_pes_22_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_28_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_28_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_28_io_in_stage = local_pes_23_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_29_clock = clock;
  assign local_pes_23_29_reset = reset;
  assign local_pes_23_29_io_in_q = local_pes_23_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_29_io_in_sum = local_pes_23_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_29_io_in_sum_exp = local_pes_23_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_29_io_in_kv = local_pes_22_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_29_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_29_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_29_io_in_stage = local_pes_23_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_30_clock = clock;
  assign local_pes_23_30_reset = reset;
  assign local_pes_23_30_io_in_q = local_pes_23_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_30_io_in_sum = local_pes_23_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_30_io_in_sum_exp = local_pes_23_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_30_io_in_kv = local_pes_22_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_30_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_30_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_30_io_in_stage = local_pes_23_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_23_31_clock = clock;
  assign local_pes_23_31_reset = reset;
  assign local_pes_23_31_io_in_q = local_pes_23_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_23_31_io_in_sum = local_pes_23_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_23_31_io_in_sum_exp = local_pes_23_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_23_31_io_in_kv = local_pes_22_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_23_31_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_23_31_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_23_31_io_in_stage = local_pes_23_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_0_clock = clock;
  assign local_pes_24_0_reset = reset;
  assign local_pes_24_0_io_in_q = io_q_ports_24; // @[PEArray.scala 51:37]
  assign local_pes_24_0_io_in_kv = io_kv_ports_55; // @[PEArray.scala 40:34]
  assign local_pes_24_0_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_0_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_0_io_in_stage = io_stage_ports_24; // @[PEArray.scala 52:41]
  assign local_pes_24_1_clock = clock;
  assign local_pes_24_1_reset = reset;
  assign local_pes_24_1_io_in_q = local_pes_24_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_1_io_in_sum = local_pes_24_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_24_1_io_in_kv = local_pes_23_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_1_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_1_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_1_io_in_stage = local_pes_24_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_2_clock = clock;
  assign local_pes_24_2_reset = reset;
  assign local_pes_24_2_io_in_q = local_pes_24_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_2_io_in_sum = local_pes_24_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_2_io_in_sum_exp = local_pes_24_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_2_io_in_kv = local_pes_23_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_2_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_2_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_2_io_in_stage = local_pes_24_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_3_clock = clock;
  assign local_pes_24_3_reset = reset;
  assign local_pes_24_3_io_in_q = local_pes_24_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_3_io_in_sum = local_pes_24_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_3_io_in_sum_exp = local_pes_24_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_3_io_in_kv = local_pes_23_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_3_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_3_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_3_io_in_stage = local_pes_24_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_4_clock = clock;
  assign local_pes_24_4_reset = reset;
  assign local_pes_24_4_io_in_q = local_pes_24_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_4_io_in_sum = local_pes_24_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_4_io_in_sum_exp = local_pes_24_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_4_io_in_kv = local_pes_23_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_4_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_4_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_4_io_in_stage = local_pes_24_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_5_clock = clock;
  assign local_pes_24_5_reset = reset;
  assign local_pes_24_5_io_in_q = local_pes_24_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_5_io_in_sum = local_pes_24_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_5_io_in_sum_exp = local_pes_24_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_5_io_in_kv = local_pes_23_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_5_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_5_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_5_io_in_stage = local_pes_24_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_6_clock = clock;
  assign local_pes_24_6_reset = reset;
  assign local_pes_24_6_io_in_q = local_pes_24_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_6_io_in_sum = local_pes_24_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_6_io_in_sum_exp = local_pes_24_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_6_io_in_kv = local_pes_23_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_6_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_6_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_6_io_in_stage = local_pes_24_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_7_clock = clock;
  assign local_pes_24_7_reset = reset;
  assign local_pes_24_7_io_in_q = local_pes_24_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_7_io_in_sum = local_pes_24_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_7_io_in_sum_exp = local_pes_24_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_7_io_in_kv = local_pes_23_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_7_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_7_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_7_io_in_stage = local_pes_24_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_8_clock = clock;
  assign local_pes_24_8_reset = reset;
  assign local_pes_24_8_io_in_q = local_pes_24_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_8_io_in_sum = local_pes_24_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_8_io_in_sum_exp = local_pes_24_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_8_io_in_kv = local_pes_23_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_8_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_8_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_8_io_in_stage = local_pes_24_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_9_clock = clock;
  assign local_pes_24_9_reset = reset;
  assign local_pes_24_9_io_in_q = local_pes_24_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_9_io_in_sum = local_pes_24_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_9_io_in_sum_exp = local_pes_24_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_9_io_in_kv = local_pes_23_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_9_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_9_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_9_io_in_stage = local_pes_24_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_10_clock = clock;
  assign local_pes_24_10_reset = reset;
  assign local_pes_24_10_io_in_q = local_pes_24_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_10_io_in_sum = local_pes_24_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_10_io_in_sum_exp = local_pes_24_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_10_io_in_kv = local_pes_23_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_10_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_10_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_10_io_in_stage = local_pes_24_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_11_clock = clock;
  assign local_pes_24_11_reset = reset;
  assign local_pes_24_11_io_in_q = local_pes_24_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_11_io_in_sum = local_pes_24_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_11_io_in_sum_exp = local_pes_24_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_11_io_in_kv = local_pes_23_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_11_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_11_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_11_io_in_stage = local_pes_24_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_12_clock = clock;
  assign local_pes_24_12_reset = reset;
  assign local_pes_24_12_io_in_q = local_pes_24_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_12_io_in_sum = local_pes_24_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_12_io_in_sum_exp = local_pes_24_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_12_io_in_kv = local_pes_23_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_12_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_12_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_12_io_in_stage = local_pes_24_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_13_clock = clock;
  assign local_pes_24_13_reset = reset;
  assign local_pes_24_13_io_in_q = local_pes_24_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_13_io_in_sum = local_pes_24_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_13_io_in_sum_exp = local_pes_24_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_13_io_in_kv = local_pes_23_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_13_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_13_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_13_io_in_stage = local_pes_24_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_14_clock = clock;
  assign local_pes_24_14_reset = reset;
  assign local_pes_24_14_io_in_q = local_pes_24_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_14_io_in_sum = local_pes_24_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_14_io_in_sum_exp = local_pes_24_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_14_io_in_kv = local_pes_23_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_14_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_14_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_14_io_in_stage = local_pes_24_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_15_clock = clock;
  assign local_pes_24_15_reset = reset;
  assign local_pes_24_15_io_in_q = local_pes_24_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_15_io_in_sum = local_pes_24_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_15_io_in_sum_exp = local_pes_24_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_15_io_in_kv = local_pes_23_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_15_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_15_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_15_io_in_stage = local_pes_24_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_16_clock = clock;
  assign local_pes_24_16_reset = reset;
  assign local_pes_24_16_io_in_q = local_pes_24_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_16_io_in_sum = local_pes_24_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_16_io_in_sum_exp = local_pes_24_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_16_io_in_kv = local_pes_23_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_16_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_16_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_16_io_in_stage = local_pes_24_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_17_clock = clock;
  assign local_pes_24_17_reset = reset;
  assign local_pes_24_17_io_in_q = local_pes_24_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_17_io_in_sum = local_pes_24_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_17_io_in_sum_exp = local_pes_24_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_17_io_in_kv = local_pes_23_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_17_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_17_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_17_io_in_stage = local_pes_24_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_18_clock = clock;
  assign local_pes_24_18_reset = reset;
  assign local_pes_24_18_io_in_q = local_pes_24_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_18_io_in_sum = local_pes_24_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_18_io_in_sum_exp = local_pes_24_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_18_io_in_kv = local_pes_23_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_18_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_18_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_18_io_in_stage = local_pes_24_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_19_clock = clock;
  assign local_pes_24_19_reset = reset;
  assign local_pes_24_19_io_in_q = local_pes_24_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_19_io_in_sum = local_pes_24_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_19_io_in_sum_exp = local_pes_24_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_19_io_in_kv = local_pes_23_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_19_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_19_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_19_io_in_stage = local_pes_24_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_20_clock = clock;
  assign local_pes_24_20_reset = reset;
  assign local_pes_24_20_io_in_q = local_pes_24_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_20_io_in_sum = local_pes_24_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_20_io_in_sum_exp = local_pes_24_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_20_io_in_kv = local_pes_23_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_20_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_20_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_20_io_in_stage = local_pes_24_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_21_clock = clock;
  assign local_pes_24_21_reset = reset;
  assign local_pes_24_21_io_in_q = local_pes_24_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_21_io_in_sum = local_pes_24_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_21_io_in_sum_exp = local_pes_24_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_21_io_in_kv = local_pes_23_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_21_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_21_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_21_io_in_stage = local_pes_24_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_22_clock = clock;
  assign local_pes_24_22_reset = reset;
  assign local_pes_24_22_io_in_q = local_pes_24_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_22_io_in_sum = local_pes_24_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_22_io_in_sum_exp = local_pes_24_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_22_io_in_kv = local_pes_23_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_22_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_22_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_22_io_in_stage = local_pes_24_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_23_clock = clock;
  assign local_pes_24_23_reset = reset;
  assign local_pes_24_23_io_in_q = local_pes_24_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_23_io_in_sum = local_pes_24_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_23_io_in_sum_exp = local_pes_24_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_23_io_in_kv = local_pes_23_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_23_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_23_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_23_io_in_stage = local_pes_24_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_24_clock = clock;
  assign local_pes_24_24_reset = reset;
  assign local_pes_24_24_io_in_q = local_pes_24_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_24_io_in_sum = local_pes_24_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_24_io_in_sum_exp = local_pes_24_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_24_io_in_kv = local_pes_23_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_24_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_24_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_24_io_in_stage = local_pes_24_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_25_clock = clock;
  assign local_pes_24_25_reset = reset;
  assign local_pes_24_25_io_in_q = local_pes_24_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_25_io_in_sum = local_pes_24_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_25_io_in_sum_exp = local_pes_24_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_25_io_in_kv = local_pes_23_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_25_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_25_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_25_io_in_stage = local_pes_24_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_26_clock = clock;
  assign local_pes_24_26_reset = reset;
  assign local_pes_24_26_io_in_q = local_pes_24_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_26_io_in_sum = local_pes_24_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_26_io_in_sum_exp = local_pes_24_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_26_io_in_kv = local_pes_23_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_26_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_26_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_26_io_in_stage = local_pes_24_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_27_clock = clock;
  assign local_pes_24_27_reset = reset;
  assign local_pes_24_27_io_in_q = local_pes_24_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_27_io_in_sum = local_pes_24_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_27_io_in_sum_exp = local_pes_24_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_27_io_in_kv = local_pes_23_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_27_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_27_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_27_io_in_stage = local_pes_24_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_28_clock = clock;
  assign local_pes_24_28_reset = reset;
  assign local_pes_24_28_io_in_q = local_pes_24_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_28_io_in_sum = local_pes_24_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_28_io_in_sum_exp = local_pes_24_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_28_io_in_kv = local_pes_23_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_28_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_28_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_28_io_in_stage = local_pes_24_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_29_clock = clock;
  assign local_pes_24_29_reset = reset;
  assign local_pes_24_29_io_in_q = local_pes_24_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_29_io_in_sum = local_pes_24_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_29_io_in_sum_exp = local_pes_24_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_29_io_in_kv = local_pes_23_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_29_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_29_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_29_io_in_stage = local_pes_24_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_30_clock = clock;
  assign local_pes_24_30_reset = reset;
  assign local_pes_24_30_io_in_q = local_pes_24_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_30_io_in_sum = local_pes_24_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_30_io_in_sum_exp = local_pes_24_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_30_io_in_kv = local_pes_23_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_30_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_30_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_30_io_in_stage = local_pes_24_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_24_31_clock = clock;
  assign local_pes_24_31_reset = reset;
  assign local_pes_24_31_io_in_q = local_pes_24_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_24_31_io_in_sum = local_pes_24_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_24_31_io_in_sum_exp = local_pes_24_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_24_31_io_in_kv = local_pes_23_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_24_31_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_24_31_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_24_31_io_in_stage = local_pes_24_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_0_clock = clock;
  assign local_pes_25_0_reset = reset;
  assign local_pes_25_0_io_in_q = io_q_ports_25; // @[PEArray.scala 51:37]
  assign local_pes_25_0_io_in_kv = io_kv_ports_56; // @[PEArray.scala 40:34]
  assign local_pes_25_0_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_0_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_0_io_in_stage = io_stage_ports_25; // @[PEArray.scala 52:41]
  assign local_pes_25_1_clock = clock;
  assign local_pes_25_1_reset = reset;
  assign local_pes_25_1_io_in_q = local_pes_25_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_1_io_in_sum = local_pes_25_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_25_1_io_in_kv = local_pes_24_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_1_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_1_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_1_io_in_stage = local_pes_25_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_2_clock = clock;
  assign local_pes_25_2_reset = reset;
  assign local_pes_25_2_io_in_q = local_pes_25_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_2_io_in_sum = local_pes_25_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_2_io_in_sum_exp = local_pes_25_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_2_io_in_kv = local_pes_24_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_2_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_2_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_2_io_in_stage = local_pes_25_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_3_clock = clock;
  assign local_pes_25_3_reset = reset;
  assign local_pes_25_3_io_in_q = local_pes_25_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_3_io_in_sum = local_pes_25_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_3_io_in_sum_exp = local_pes_25_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_3_io_in_kv = local_pes_24_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_3_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_3_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_3_io_in_stage = local_pes_25_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_4_clock = clock;
  assign local_pes_25_4_reset = reset;
  assign local_pes_25_4_io_in_q = local_pes_25_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_4_io_in_sum = local_pes_25_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_4_io_in_sum_exp = local_pes_25_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_4_io_in_kv = local_pes_24_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_4_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_4_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_4_io_in_stage = local_pes_25_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_5_clock = clock;
  assign local_pes_25_5_reset = reset;
  assign local_pes_25_5_io_in_q = local_pes_25_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_5_io_in_sum = local_pes_25_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_5_io_in_sum_exp = local_pes_25_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_5_io_in_kv = local_pes_24_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_5_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_5_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_5_io_in_stage = local_pes_25_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_6_clock = clock;
  assign local_pes_25_6_reset = reset;
  assign local_pes_25_6_io_in_q = local_pes_25_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_6_io_in_sum = local_pes_25_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_6_io_in_sum_exp = local_pes_25_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_6_io_in_kv = local_pes_24_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_6_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_6_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_6_io_in_stage = local_pes_25_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_7_clock = clock;
  assign local_pes_25_7_reset = reset;
  assign local_pes_25_7_io_in_q = local_pes_25_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_7_io_in_sum = local_pes_25_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_7_io_in_sum_exp = local_pes_25_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_7_io_in_kv = local_pes_24_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_7_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_7_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_7_io_in_stage = local_pes_25_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_8_clock = clock;
  assign local_pes_25_8_reset = reset;
  assign local_pes_25_8_io_in_q = local_pes_25_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_8_io_in_sum = local_pes_25_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_8_io_in_sum_exp = local_pes_25_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_8_io_in_kv = local_pes_24_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_8_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_8_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_8_io_in_stage = local_pes_25_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_9_clock = clock;
  assign local_pes_25_9_reset = reset;
  assign local_pes_25_9_io_in_q = local_pes_25_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_9_io_in_sum = local_pes_25_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_9_io_in_sum_exp = local_pes_25_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_9_io_in_kv = local_pes_24_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_9_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_9_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_9_io_in_stage = local_pes_25_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_10_clock = clock;
  assign local_pes_25_10_reset = reset;
  assign local_pes_25_10_io_in_q = local_pes_25_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_10_io_in_sum = local_pes_25_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_10_io_in_sum_exp = local_pes_25_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_10_io_in_kv = local_pes_24_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_10_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_10_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_10_io_in_stage = local_pes_25_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_11_clock = clock;
  assign local_pes_25_11_reset = reset;
  assign local_pes_25_11_io_in_q = local_pes_25_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_11_io_in_sum = local_pes_25_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_11_io_in_sum_exp = local_pes_25_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_11_io_in_kv = local_pes_24_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_11_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_11_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_11_io_in_stage = local_pes_25_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_12_clock = clock;
  assign local_pes_25_12_reset = reset;
  assign local_pes_25_12_io_in_q = local_pes_25_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_12_io_in_sum = local_pes_25_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_12_io_in_sum_exp = local_pes_25_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_12_io_in_kv = local_pes_24_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_12_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_12_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_12_io_in_stage = local_pes_25_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_13_clock = clock;
  assign local_pes_25_13_reset = reset;
  assign local_pes_25_13_io_in_q = local_pes_25_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_13_io_in_sum = local_pes_25_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_13_io_in_sum_exp = local_pes_25_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_13_io_in_kv = local_pes_24_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_13_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_13_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_13_io_in_stage = local_pes_25_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_14_clock = clock;
  assign local_pes_25_14_reset = reset;
  assign local_pes_25_14_io_in_q = local_pes_25_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_14_io_in_sum = local_pes_25_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_14_io_in_sum_exp = local_pes_25_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_14_io_in_kv = local_pes_24_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_14_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_14_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_14_io_in_stage = local_pes_25_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_15_clock = clock;
  assign local_pes_25_15_reset = reset;
  assign local_pes_25_15_io_in_q = local_pes_25_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_15_io_in_sum = local_pes_25_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_15_io_in_sum_exp = local_pes_25_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_15_io_in_kv = local_pes_24_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_15_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_15_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_15_io_in_stage = local_pes_25_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_16_clock = clock;
  assign local_pes_25_16_reset = reset;
  assign local_pes_25_16_io_in_q = local_pes_25_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_16_io_in_sum = local_pes_25_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_16_io_in_sum_exp = local_pes_25_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_16_io_in_kv = local_pes_24_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_16_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_16_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_16_io_in_stage = local_pes_25_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_17_clock = clock;
  assign local_pes_25_17_reset = reset;
  assign local_pes_25_17_io_in_q = local_pes_25_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_17_io_in_sum = local_pes_25_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_17_io_in_sum_exp = local_pes_25_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_17_io_in_kv = local_pes_24_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_17_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_17_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_17_io_in_stage = local_pes_25_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_18_clock = clock;
  assign local_pes_25_18_reset = reset;
  assign local_pes_25_18_io_in_q = local_pes_25_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_18_io_in_sum = local_pes_25_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_18_io_in_sum_exp = local_pes_25_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_18_io_in_kv = local_pes_24_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_18_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_18_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_18_io_in_stage = local_pes_25_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_19_clock = clock;
  assign local_pes_25_19_reset = reset;
  assign local_pes_25_19_io_in_q = local_pes_25_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_19_io_in_sum = local_pes_25_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_19_io_in_sum_exp = local_pes_25_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_19_io_in_kv = local_pes_24_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_19_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_19_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_19_io_in_stage = local_pes_25_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_20_clock = clock;
  assign local_pes_25_20_reset = reset;
  assign local_pes_25_20_io_in_q = local_pes_25_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_20_io_in_sum = local_pes_25_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_20_io_in_sum_exp = local_pes_25_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_20_io_in_kv = local_pes_24_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_20_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_20_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_20_io_in_stage = local_pes_25_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_21_clock = clock;
  assign local_pes_25_21_reset = reset;
  assign local_pes_25_21_io_in_q = local_pes_25_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_21_io_in_sum = local_pes_25_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_21_io_in_sum_exp = local_pes_25_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_21_io_in_kv = local_pes_24_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_21_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_21_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_21_io_in_stage = local_pes_25_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_22_clock = clock;
  assign local_pes_25_22_reset = reset;
  assign local_pes_25_22_io_in_q = local_pes_25_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_22_io_in_sum = local_pes_25_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_22_io_in_sum_exp = local_pes_25_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_22_io_in_kv = local_pes_24_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_22_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_22_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_22_io_in_stage = local_pes_25_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_23_clock = clock;
  assign local_pes_25_23_reset = reset;
  assign local_pes_25_23_io_in_q = local_pes_25_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_23_io_in_sum = local_pes_25_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_23_io_in_sum_exp = local_pes_25_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_23_io_in_kv = local_pes_24_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_23_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_23_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_23_io_in_stage = local_pes_25_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_24_clock = clock;
  assign local_pes_25_24_reset = reset;
  assign local_pes_25_24_io_in_q = local_pes_25_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_24_io_in_sum = local_pes_25_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_24_io_in_sum_exp = local_pes_25_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_24_io_in_kv = local_pes_24_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_24_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_24_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_24_io_in_stage = local_pes_25_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_25_clock = clock;
  assign local_pes_25_25_reset = reset;
  assign local_pes_25_25_io_in_q = local_pes_25_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_25_io_in_sum = local_pes_25_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_25_io_in_sum_exp = local_pes_25_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_25_io_in_kv = local_pes_24_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_25_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_25_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_25_io_in_stage = local_pes_25_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_26_clock = clock;
  assign local_pes_25_26_reset = reset;
  assign local_pes_25_26_io_in_q = local_pes_25_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_26_io_in_sum = local_pes_25_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_26_io_in_sum_exp = local_pes_25_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_26_io_in_kv = local_pes_24_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_26_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_26_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_26_io_in_stage = local_pes_25_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_27_clock = clock;
  assign local_pes_25_27_reset = reset;
  assign local_pes_25_27_io_in_q = local_pes_25_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_27_io_in_sum = local_pes_25_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_27_io_in_sum_exp = local_pes_25_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_27_io_in_kv = local_pes_24_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_27_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_27_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_27_io_in_stage = local_pes_25_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_28_clock = clock;
  assign local_pes_25_28_reset = reset;
  assign local_pes_25_28_io_in_q = local_pes_25_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_28_io_in_sum = local_pes_25_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_28_io_in_sum_exp = local_pes_25_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_28_io_in_kv = local_pes_24_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_28_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_28_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_28_io_in_stage = local_pes_25_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_29_clock = clock;
  assign local_pes_25_29_reset = reset;
  assign local_pes_25_29_io_in_q = local_pes_25_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_29_io_in_sum = local_pes_25_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_29_io_in_sum_exp = local_pes_25_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_29_io_in_kv = local_pes_24_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_29_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_29_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_29_io_in_stage = local_pes_25_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_30_clock = clock;
  assign local_pes_25_30_reset = reset;
  assign local_pes_25_30_io_in_q = local_pes_25_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_30_io_in_sum = local_pes_25_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_30_io_in_sum_exp = local_pes_25_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_30_io_in_kv = local_pes_24_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_30_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_30_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_30_io_in_stage = local_pes_25_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_25_31_clock = clock;
  assign local_pes_25_31_reset = reset;
  assign local_pes_25_31_io_in_q = local_pes_25_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_25_31_io_in_sum = local_pes_25_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_25_31_io_in_sum_exp = local_pes_25_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_25_31_io_in_kv = local_pes_24_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_25_31_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_25_31_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_25_31_io_in_stage = local_pes_25_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_0_clock = clock;
  assign local_pes_26_0_reset = reset;
  assign local_pes_26_0_io_in_q = io_q_ports_26; // @[PEArray.scala 51:37]
  assign local_pes_26_0_io_in_kv = io_kv_ports_57; // @[PEArray.scala 40:34]
  assign local_pes_26_0_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_0_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_0_io_in_stage = io_stage_ports_26; // @[PEArray.scala 52:41]
  assign local_pes_26_1_clock = clock;
  assign local_pes_26_1_reset = reset;
  assign local_pes_26_1_io_in_q = local_pes_26_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_1_io_in_sum = local_pes_26_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_26_1_io_in_kv = local_pes_25_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_1_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_1_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_1_io_in_stage = local_pes_26_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_2_clock = clock;
  assign local_pes_26_2_reset = reset;
  assign local_pes_26_2_io_in_q = local_pes_26_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_2_io_in_sum = local_pes_26_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_2_io_in_sum_exp = local_pes_26_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_2_io_in_kv = local_pes_25_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_2_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_2_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_2_io_in_stage = local_pes_26_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_3_clock = clock;
  assign local_pes_26_3_reset = reset;
  assign local_pes_26_3_io_in_q = local_pes_26_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_3_io_in_sum = local_pes_26_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_3_io_in_sum_exp = local_pes_26_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_3_io_in_kv = local_pes_25_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_3_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_3_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_3_io_in_stage = local_pes_26_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_4_clock = clock;
  assign local_pes_26_4_reset = reset;
  assign local_pes_26_4_io_in_q = local_pes_26_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_4_io_in_sum = local_pes_26_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_4_io_in_sum_exp = local_pes_26_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_4_io_in_kv = local_pes_25_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_4_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_4_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_4_io_in_stage = local_pes_26_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_5_clock = clock;
  assign local_pes_26_5_reset = reset;
  assign local_pes_26_5_io_in_q = local_pes_26_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_5_io_in_sum = local_pes_26_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_5_io_in_sum_exp = local_pes_26_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_5_io_in_kv = local_pes_25_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_5_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_5_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_5_io_in_stage = local_pes_26_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_6_clock = clock;
  assign local_pes_26_6_reset = reset;
  assign local_pes_26_6_io_in_q = local_pes_26_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_6_io_in_sum = local_pes_26_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_6_io_in_sum_exp = local_pes_26_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_6_io_in_kv = local_pes_25_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_6_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_6_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_6_io_in_stage = local_pes_26_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_7_clock = clock;
  assign local_pes_26_7_reset = reset;
  assign local_pes_26_7_io_in_q = local_pes_26_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_7_io_in_sum = local_pes_26_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_7_io_in_sum_exp = local_pes_26_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_7_io_in_kv = local_pes_25_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_7_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_7_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_7_io_in_stage = local_pes_26_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_8_clock = clock;
  assign local_pes_26_8_reset = reset;
  assign local_pes_26_8_io_in_q = local_pes_26_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_8_io_in_sum = local_pes_26_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_8_io_in_sum_exp = local_pes_26_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_8_io_in_kv = local_pes_25_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_8_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_8_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_8_io_in_stage = local_pes_26_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_9_clock = clock;
  assign local_pes_26_9_reset = reset;
  assign local_pes_26_9_io_in_q = local_pes_26_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_9_io_in_sum = local_pes_26_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_9_io_in_sum_exp = local_pes_26_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_9_io_in_kv = local_pes_25_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_9_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_9_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_9_io_in_stage = local_pes_26_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_10_clock = clock;
  assign local_pes_26_10_reset = reset;
  assign local_pes_26_10_io_in_q = local_pes_26_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_10_io_in_sum = local_pes_26_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_10_io_in_sum_exp = local_pes_26_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_10_io_in_kv = local_pes_25_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_10_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_10_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_10_io_in_stage = local_pes_26_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_11_clock = clock;
  assign local_pes_26_11_reset = reset;
  assign local_pes_26_11_io_in_q = local_pes_26_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_11_io_in_sum = local_pes_26_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_11_io_in_sum_exp = local_pes_26_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_11_io_in_kv = local_pes_25_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_11_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_11_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_11_io_in_stage = local_pes_26_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_12_clock = clock;
  assign local_pes_26_12_reset = reset;
  assign local_pes_26_12_io_in_q = local_pes_26_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_12_io_in_sum = local_pes_26_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_12_io_in_sum_exp = local_pes_26_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_12_io_in_kv = local_pes_25_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_12_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_12_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_12_io_in_stage = local_pes_26_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_13_clock = clock;
  assign local_pes_26_13_reset = reset;
  assign local_pes_26_13_io_in_q = local_pes_26_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_13_io_in_sum = local_pes_26_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_13_io_in_sum_exp = local_pes_26_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_13_io_in_kv = local_pes_25_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_13_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_13_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_13_io_in_stage = local_pes_26_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_14_clock = clock;
  assign local_pes_26_14_reset = reset;
  assign local_pes_26_14_io_in_q = local_pes_26_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_14_io_in_sum = local_pes_26_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_14_io_in_sum_exp = local_pes_26_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_14_io_in_kv = local_pes_25_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_14_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_14_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_14_io_in_stage = local_pes_26_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_15_clock = clock;
  assign local_pes_26_15_reset = reset;
  assign local_pes_26_15_io_in_q = local_pes_26_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_15_io_in_sum = local_pes_26_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_15_io_in_sum_exp = local_pes_26_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_15_io_in_kv = local_pes_25_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_15_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_15_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_15_io_in_stage = local_pes_26_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_16_clock = clock;
  assign local_pes_26_16_reset = reset;
  assign local_pes_26_16_io_in_q = local_pes_26_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_16_io_in_sum = local_pes_26_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_16_io_in_sum_exp = local_pes_26_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_16_io_in_kv = local_pes_25_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_16_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_16_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_16_io_in_stage = local_pes_26_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_17_clock = clock;
  assign local_pes_26_17_reset = reset;
  assign local_pes_26_17_io_in_q = local_pes_26_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_17_io_in_sum = local_pes_26_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_17_io_in_sum_exp = local_pes_26_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_17_io_in_kv = local_pes_25_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_17_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_17_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_17_io_in_stage = local_pes_26_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_18_clock = clock;
  assign local_pes_26_18_reset = reset;
  assign local_pes_26_18_io_in_q = local_pes_26_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_18_io_in_sum = local_pes_26_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_18_io_in_sum_exp = local_pes_26_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_18_io_in_kv = local_pes_25_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_18_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_18_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_18_io_in_stage = local_pes_26_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_19_clock = clock;
  assign local_pes_26_19_reset = reset;
  assign local_pes_26_19_io_in_q = local_pes_26_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_19_io_in_sum = local_pes_26_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_19_io_in_sum_exp = local_pes_26_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_19_io_in_kv = local_pes_25_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_19_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_19_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_19_io_in_stage = local_pes_26_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_20_clock = clock;
  assign local_pes_26_20_reset = reset;
  assign local_pes_26_20_io_in_q = local_pes_26_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_20_io_in_sum = local_pes_26_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_20_io_in_sum_exp = local_pes_26_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_20_io_in_kv = local_pes_25_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_20_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_20_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_20_io_in_stage = local_pes_26_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_21_clock = clock;
  assign local_pes_26_21_reset = reset;
  assign local_pes_26_21_io_in_q = local_pes_26_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_21_io_in_sum = local_pes_26_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_21_io_in_sum_exp = local_pes_26_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_21_io_in_kv = local_pes_25_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_21_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_21_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_21_io_in_stage = local_pes_26_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_22_clock = clock;
  assign local_pes_26_22_reset = reset;
  assign local_pes_26_22_io_in_q = local_pes_26_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_22_io_in_sum = local_pes_26_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_22_io_in_sum_exp = local_pes_26_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_22_io_in_kv = local_pes_25_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_22_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_22_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_22_io_in_stage = local_pes_26_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_23_clock = clock;
  assign local_pes_26_23_reset = reset;
  assign local_pes_26_23_io_in_q = local_pes_26_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_23_io_in_sum = local_pes_26_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_23_io_in_sum_exp = local_pes_26_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_23_io_in_kv = local_pes_25_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_23_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_23_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_23_io_in_stage = local_pes_26_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_24_clock = clock;
  assign local_pes_26_24_reset = reset;
  assign local_pes_26_24_io_in_q = local_pes_26_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_24_io_in_sum = local_pes_26_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_24_io_in_sum_exp = local_pes_26_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_24_io_in_kv = local_pes_25_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_24_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_24_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_24_io_in_stage = local_pes_26_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_25_clock = clock;
  assign local_pes_26_25_reset = reset;
  assign local_pes_26_25_io_in_q = local_pes_26_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_25_io_in_sum = local_pes_26_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_25_io_in_sum_exp = local_pes_26_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_25_io_in_kv = local_pes_25_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_25_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_25_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_25_io_in_stage = local_pes_26_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_26_clock = clock;
  assign local_pes_26_26_reset = reset;
  assign local_pes_26_26_io_in_q = local_pes_26_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_26_io_in_sum = local_pes_26_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_26_io_in_sum_exp = local_pes_26_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_26_io_in_kv = local_pes_25_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_26_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_26_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_26_io_in_stage = local_pes_26_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_27_clock = clock;
  assign local_pes_26_27_reset = reset;
  assign local_pes_26_27_io_in_q = local_pes_26_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_27_io_in_sum = local_pes_26_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_27_io_in_sum_exp = local_pes_26_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_27_io_in_kv = local_pes_25_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_27_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_27_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_27_io_in_stage = local_pes_26_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_28_clock = clock;
  assign local_pes_26_28_reset = reset;
  assign local_pes_26_28_io_in_q = local_pes_26_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_28_io_in_sum = local_pes_26_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_28_io_in_sum_exp = local_pes_26_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_28_io_in_kv = local_pes_25_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_28_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_28_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_28_io_in_stage = local_pes_26_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_29_clock = clock;
  assign local_pes_26_29_reset = reset;
  assign local_pes_26_29_io_in_q = local_pes_26_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_29_io_in_sum = local_pes_26_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_29_io_in_sum_exp = local_pes_26_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_29_io_in_kv = local_pes_25_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_29_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_29_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_29_io_in_stage = local_pes_26_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_30_clock = clock;
  assign local_pes_26_30_reset = reset;
  assign local_pes_26_30_io_in_q = local_pes_26_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_30_io_in_sum = local_pes_26_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_30_io_in_sum_exp = local_pes_26_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_30_io_in_kv = local_pes_25_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_30_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_30_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_30_io_in_stage = local_pes_26_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_26_31_clock = clock;
  assign local_pes_26_31_reset = reset;
  assign local_pes_26_31_io_in_q = local_pes_26_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_26_31_io_in_sum = local_pes_26_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_26_31_io_in_sum_exp = local_pes_26_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_26_31_io_in_kv = local_pes_25_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_26_31_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_26_31_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_26_31_io_in_stage = local_pes_26_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_0_clock = clock;
  assign local_pes_27_0_reset = reset;
  assign local_pes_27_0_io_in_q = io_q_ports_27; // @[PEArray.scala 51:37]
  assign local_pes_27_0_io_in_kv = io_kv_ports_58; // @[PEArray.scala 40:34]
  assign local_pes_27_0_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_0_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_0_io_in_stage = io_stage_ports_27; // @[PEArray.scala 52:41]
  assign local_pes_27_1_clock = clock;
  assign local_pes_27_1_reset = reset;
  assign local_pes_27_1_io_in_q = local_pes_27_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_1_io_in_sum = local_pes_27_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_27_1_io_in_kv = local_pes_26_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_1_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_1_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_1_io_in_stage = local_pes_27_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_2_clock = clock;
  assign local_pes_27_2_reset = reset;
  assign local_pes_27_2_io_in_q = local_pes_27_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_2_io_in_sum = local_pes_27_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_2_io_in_sum_exp = local_pes_27_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_2_io_in_kv = local_pes_26_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_2_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_2_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_2_io_in_stage = local_pes_27_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_3_clock = clock;
  assign local_pes_27_3_reset = reset;
  assign local_pes_27_3_io_in_q = local_pes_27_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_3_io_in_sum = local_pes_27_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_3_io_in_sum_exp = local_pes_27_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_3_io_in_kv = local_pes_26_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_3_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_3_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_3_io_in_stage = local_pes_27_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_4_clock = clock;
  assign local_pes_27_4_reset = reset;
  assign local_pes_27_4_io_in_q = local_pes_27_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_4_io_in_sum = local_pes_27_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_4_io_in_sum_exp = local_pes_27_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_4_io_in_kv = local_pes_26_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_4_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_4_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_4_io_in_stage = local_pes_27_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_5_clock = clock;
  assign local_pes_27_5_reset = reset;
  assign local_pes_27_5_io_in_q = local_pes_27_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_5_io_in_sum = local_pes_27_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_5_io_in_sum_exp = local_pes_27_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_5_io_in_kv = local_pes_26_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_5_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_5_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_5_io_in_stage = local_pes_27_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_6_clock = clock;
  assign local_pes_27_6_reset = reset;
  assign local_pes_27_6_io_in_q = local_pes_27_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_6_io_in_sum = local_pes_27_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_6_io_in_sum_exp = local_pes_27_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_6_io_in_kv = local_pes_26_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_6_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_6_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_6_io_in_stage = local_pes_27_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_7_clock = clock;
  assign local_pes_27_7_reset = reset;
  assign local_pes_27_7_io_in_q = local_pes_27_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_7_io_in_sum = local_pes_27_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_7_io_in_sum_exp = local_pes_27_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_7_io_in_kv = local_pes_26_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_7_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_7_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_7_io_in_stage = local_pes_27_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_8_clock = clock;
  assign local_pes_27_8_reset = reset;
  assign local_pes_27_8_io_in_q = local_pes_27_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_8_io_in_sum = local_pes_27_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_8_io_in_sum_exp = local_pes_27_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_8_io_in_kv = local_pes_26_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_8_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_8_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_8_io_in_stage = local_pes_27_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_9_clock = clock;
  assign local_pes_27_9_reset = reset;
  assign local_pes_27_9_io_in_q = local_pes_27_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_9_io_in_sum = local_pes_27_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_9_io_in_sum_exp = local_pes_27_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_9_io_in_kv = local_pes_26_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_9_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_9_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_9_io_in_stage = local_pes_27_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_10_clock = clock;
  assign local_pes_27_10_reset = reset;
  assign local_pes_27_10_io_in_q = local_pes_27_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_10_io_in_sum = local_pes_27_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_10_io_in_sum_exp = local_pes_27_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_10_io_in_kv = local_pes_26_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_10_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_10_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_10_io_in_stage = local_pes_27_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_11_clock = clock;
  assign local_pes_27_11_reset = reset;
  assign local_pes_27_11_io_in_q = local_pes_27_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_11_io_in_sum = local_pes_27_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_11_io_in_sum_exp = local_pes_27_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_11_io_in_kv = local_pes_26_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_11_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_11_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_11_io_in_stage = local_pes_27_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_12_clock = clock;
  assign local_pes_27_12_reset = reset;
  assign local_pes_27_12_io_in_q = local_pes_27_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_12_io_in_sum = local_pes_27_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_12_io_in_sum_exp = local_pes_27_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_12_io_in_kv = local_pes_26_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_12_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_12_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_12_io_in_stage = local_pes_27_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_13_clock = clock;
  assign local_pes_27_13_reset = reset;
  assign local_pes_27_13_io_in_q = local_pes_27_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_13_io_in_sum = local_pes_27_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_13_io_in_sum_exp = local_pes_27_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_13_io_in_kv = local_pes_26_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_13_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_13_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_13_io_in_stage = local_pes_27_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_14_clock = clock;
  assign local_pes_27_14_reset = reset;
  assign local_pes_27_14_io_in_q = local_pes_27_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_14_io_in_sum = local_pes_27_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_14_io_in_sum_exp = local_pes_27_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_14_io_in_kv = local_pes_26_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_14_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_14_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_14_io_in_stage = local_pes_27_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_15_clock = clock;
  assign local_pes_27_15_reset = reset;
  assign local_pes_27_15_io_in_q = local_pes_27_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_15_io_in_sum = local_pes_27_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_15_io_in_sum_exp = local_pes_27_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_15_io_in_kv = local_pes_26_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_15_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_15_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_15_io_in_stage = local_pes_27_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_16_clock = clock;
  assign local_pes_27_16_reset = reset;
  assign local_pes_27_16_io_in_q = local_pes_27_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_16_io_in_sum = local_pes_27_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_16_io_in_sum_exp = local_pes_27_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_16_io_in_kv = local_pes_26_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_16_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_16_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_16_io_in_stage = local_pes_27_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_17_clock = clock;
  assign local_pes_27_17_reset = reset;
  assign local_pes_27_17_io_in_q = local_pes_27_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_17_io_in_sum = local_pes_27_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_17_io_in_sum_exp = local_pes_27_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_17_io_in_kv = local_pes_26_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_17_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_17_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_17_io_in_stage = local_pes_27_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_18_clock = clock;
  assign local_pes_27_18_reset = reset;
  assign local_pes_27_18_io_in_q = local_pes_27_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_18_io_in_sum = local_pes_27_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_18_io_in_sum_exp = local_pes_27_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_18_io_in_kv = local_pes_26_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_18_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_18_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_18_io_in_stage = local_pes_27_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_19_clock = clock;
  assign local_pes_27_19_reset = reset;
  assign local_pes_27_19_io_in_q = local_pes_27_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_19_io_in_sum = local_pes_27_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_19_io_in_sum_exp = local_pes_27_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_19_io_in_kv = local_pes_26_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_19_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_19_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_19_io_in_stage = local_pes_27_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_20_clock = clock;
  assign local_pes_27_20_reset = reset;
  assign local_pes_27_20_io_in_q = local_pes_27_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_20_io_in_sum = local_pes_27_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_20_io_in_sum_exp = local_pes_27_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_20_io_in_kv = local_pes_26_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_20_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_20_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_20_io_in_stage = local_pes_27_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_21_clock = clock;
  assign local_pes_27_21_reset = reset;
  assign local_pes_27_21_io_in_q = local_pes_27_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_21_io_in_sum = local_pes_27_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_21_io_in_sum_exp = local_pes_27_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_21_io_in_kv = local_pes_26_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_21_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_21_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_21_io_in_stage = local_pes_27_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_22_clock = clock;
  assign local_pes_27_22_reset = reset;
  assign local_pes_27_22_io_in_q = local_pes_27_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_22_io_in_sum = local_pes_27_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_22_io_in_sum_exp = local_pes_27_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_22_io_in_kv = local_pes_26_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_22_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_22_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_22_io_in_stage = local_pes_27_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_23_clock = clock;
  assign local_pes_27_23_reset = reset;
  assign local_pes_27_23_io_in_q = local_pes_27_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_23_io_in_sum = local_pes_27_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_23_io_in_sum_exp = local_pes_27_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_23_io_in_kv = local_pes_26_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_23_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_23_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_23_io_in_stage = local_pes_27_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_24_clock = clock;
  assign local_pes_27_24_reset = reset;
  assign local_pes_27_24_io_in_q = local_pes_27_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_24_io_in_sum = local_pes_27_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_24_io_in_sum_exp = local_pes_27_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_24_io_in_kv = local_pes_26_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_24_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_24_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_24_io_in_stage = local_pes_27_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_25_clock = clock;
  assign local_pes_27_25_reset = reset;
  assign local_pes_27_25_io_in_q = local_pes_27_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_25_io_in_sum = local_pes_27_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_25_io_in_sum_exp = local_pes_27_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_25_io_in_kv = local_pes_26_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_25_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_25_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_25_io_in_stage = local_pes_27_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_26_clock = clock;
  assign local_pes_27_26_reset = reset;
  assign local_pes_27_26_io_in_q = local_pes_27_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_26_io_in_sum = local_pes_27_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_26_io_in_sum_exp = local_pes_27_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_26_io_in_kv = local_pes_26_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_26_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_26_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_26_io_in_stage = local_pes_27_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_27_clock = clock;
  assign local_pes_27_27_reset = reset;
  assign local_pes_27_27_io_in_q = local_pes_27_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_27_io_in_sum = local_pes_27_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_27_io_in_sum_exp = local_pes_27_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_27_io_in_kv = local_pes_26_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_27_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_27_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_27_io_in_stage = local_pes_27_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_28_clock = clock;
  assign local_pes_27_28_reset = reset;
  assign local_pes_27_28_io_in_q = local_pes_27_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_28_io_in_sum = local_pes_27_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_28_io_in_sum_exp = local_pes_27_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_28_io_in_kv = local_pes_26_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_28_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_28_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_28_io_in_stage = local_pes_27_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_29_clock = clock;
  assign local_pes_27_29_reset = reset;
  assign local_pes_27_29_io_in_q = local_pes_27_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_29_io_in_sum = local_pes_27_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_29_io_in_sum_exp = local_pes_27_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_29_io_in_kv = local_pes_26_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_29_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_29_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_29_io_in_stage = local_pes_27_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_30_clock = clock;
  assign local_pes_27_30_reset = reset;
  assign local_pes_27_30_io_in_q = local_pes_27_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_30_io_in_sum = local_pes_27_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_30_io_in_sum_exp = local_pes_27_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_30_io_in_kv = local_pes_26_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_30_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_30_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_30_io_in_stage = local_pes_27_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_27_31_clock = clock;
  assign local_pes_27_31_reset = reset;
  assign local_pes_27_31_io_in_q = local_pes_27_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_27_31_io_in_sum = local_pes_27_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_27_31_io_in_sum_exp = local_pes_27_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_27_31_io_in_kv = local_pes_26_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_27_31_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_27_31_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_27_31_io_in_stage = local_pes_27_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_0_clock = clock;
  assign local_pes_28_0_reset = reset;
  assign local_pes_28_0_io_in_q = io_q_ports_28; // @[PEArray.scala 51:37]
  assign local_pes_28_0_io_in_kv = io_kv_ports_59; // @[PEArray.scala 40:34]
  assign local_pes_28_0_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_0_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_0_io_in_stage = io_stage_ports_28; // @[PEArray.scala 52:41]
  assign local_pes_28_1_clock = clock;
  assign local_pes_28_1_reset = reset;
  assign local_pes_28_1_io_in_q = local_pes_28_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_1_io_in_sum = local_pes_28_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_28_1_io_in_kv = local_pes_27_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_1_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_1_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_1_io_in_stage = local_pes_28_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_2_clock = clock;
  assign local_pes_28_2_reset = reset;
  assign local_pes_28_2_io_in_q = local_pes_28_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_2_io_in_sum = local_pes_28_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_2_io_in_sum_exp = local_pes_28_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_2_io_in_kv = local_pes_27_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_2_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_2_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_2_io_in_stage = local_pes_28_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_3_clock = clock;
  assign local_pes_28_3_reset = reset;
  assign local_pes_28_3_io_in_q = local_pes_28_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_3_io_in_sum = local_pes_28_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_3_io_in_sum_exp = local_pes_28_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_3_io_in_kv = local_pes_27_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_3_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_3_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_3_io_in_stage = local_pes_28_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_4_clock = clock;
  assign local_pes_28_4_reset = reset;
  assign local_pes_28_4_io_in_q = local_pes_28_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_4_io_in_sum = local_pes_28_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_4_io_in_sum_exp = local_pes_28_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_4_io_in_kv = local_pes_27_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_4_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_4_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_4_io_in_stage = local_pes_28_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_5_clock = clock;
  assign local_pes_28_5_reset = reset;
  assign local_pes_28_5_io_in_q = local_pes_28_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_5_io_in_sum = local_pes_28_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_5_io_in_sum_exp = local_pes_28_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_5_io_in_kv = local_pes_27_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_5_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_5_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_5_io_in_stage = local_pes_28_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_6_clock = clock;
  assign local_pes_28_6_reset = reset;
  assign local_pes_28_6_io_in_q = local_pes_28_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_6_io_in_sum = local_pes_28_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_6_io_in_sum_exp = local_pes_28_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_6_io_in_kv = local_pes_27_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_6_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_6_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_6_io_in_stage = local_pes_28_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_7_clock = clock;
  assign local_pes_28_7_reset = reset;
  assign local_pes_28_7_io_in_q = local_pes_28_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_7_io_in_sum = local_pes_28_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_7_io_in_sum_exp = local_pes_28_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_7_io_in_kv = local_pes_27_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_7_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_7_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_7_io_in_stage = local_pes_28_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_8_clock = clock;
  assign local_pes_28_8_reset = reset;
  assign local_pes_28_8_io_in_q = local_pes_28_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_8_io_in_sum = local_pes_28_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_8_io_in_sum_exp = local_pes_28_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_8_io_in_kv = local_pes_27_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_8_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_8_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_8_io_in_stage = local_pes_28_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_9_clock = clock;
  assign local_pes_28_9_reset = reset;
  assign local_pes_28_9_io_in_q = local_pes_28_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_9_io_in_sum = local_pes_28_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_9_io_in_sum_exp = local_pes_28_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_9_io_in_kv = local_pes_27_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_9_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_9_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_9_io_in_stage = local_pes_28_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_10_clock = clock;
  assign local_pes_28_10_reset = reset;
  assign local_pes_28_10_io_in_q = local_pes_28_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_10_io_in_sum = local_pes_28_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_10_io_in_sum_exp = local_pes_28_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_10_io_in_kv = local_pes_27_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_10_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_10_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_10_io_in_stage = local_pes_28_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_11_clock = clock;
  assign local_pes_28_11_reset = reset;
  assign local_pes_28_11_io_in_q = local_pes_28_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_11_io_in_sum = local_pes_28_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_11_io_in_sum_exp = local_pes_28_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_11_io_in_kv = local_pes_27_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_11_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_11_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_11_io_in_stage = local_pes_28_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_12_clock = clock;
  assign local_pes_28_12_reset = reset;
  assign local_pes_28_12_io_in_q = local_pes_28_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_12_io_in_sum = local_pes_28_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_12_io_in_sum_exp = local_pes_28_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_12_io_in_kv = local_pes_27_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_12_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_12_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_12_io_in_stage = local_pes_28_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_13_clock = clock;
  assign local_pes_28_13_reset = reset;
  assign local_pes_28_13_io_in_q = local_pes_28_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_13_io_in_sum = local_pes_28_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_13_io_in_sum_exp = local_pes_28_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_13_io_in_kv = local_pes_27_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_13_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_13_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_13_io_in_stage = local_pes_28_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_14_clock = clock;
  assign local_pes_28_14_reset = reset;
  assign local_pes_28_14_io_in_q = local_pes_28_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_14_io_in_sum = local_pes_28_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_14_io_in_sum_exp = local_pes_28_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_14_io_in_kv = local_pes_27_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_14_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_14_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_14_io_in_stage = local_pes_28_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_15_clock = clock;
  assign local_pes_28_15_reset = reset;
  assign local_pes_28_15_io_in_q = local_pes_28_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_15_io_in_sum = local_pes_28_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_15_io_in_sum_exp = local_pes_28_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_15_io_in_kv = local_pes_27_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_15_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_15_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_15_io_in_stage = local_pes_28_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_16_clock = clock;
  assign local_pes_28_16_reset = reset;
  assign local_pes_28_16_io_in_q = local_pes_28_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_16_io_in_sum = local_pes_28_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_16_io_in_sum_exp = local_pes_28_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_16_io_in_kv = local_pes_27_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_16_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_16_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_16_io_in_stage = local_pes_28_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_17_clock = clock;
  assign local_pes_28_17_reset = reset;
  assign local_pes_28_17_io_in_q = local_pes_28_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_17_io_in_sum = local_pes_28_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_17_io_in_sum_exp = local_pes_28_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_17_io_in_kv = local_pes_27_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_17_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_17_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_17_io_in_stage = local_pes_28_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_18_clock = clock;
  assign local_pes_28_18_reset = reset;
  assign local_pes_28_18_io_in_q = local_pes_28_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_18_io_in_sum = local_pes_28_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_18_io_in_sum_exp = local_pes_28_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_18_io_in_kv = local_pes_27_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_18_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_18_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_18_io_in_stage = local_pes_28_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_19_clock = clock;
  assign local_pes_28_19_reset = reset;
  assign local_pes_28_19_io_in_q = local_pes_28_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_19_io_in_sum = local_pes_28_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_19_io_in_sum_exp = local_pes_28_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_19_io_in_kv = local_pes_27_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_19_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_19_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_19_io_in_stage = local_pes_28_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_20_clock = clock;
  assign local_pes_28_20_reset = reset;
  assign local_pes_28_20_io_in_q = local_pes_28_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_20_io_in_sum = local_pes_28_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_20_io_in_sum_exp = local_pes_28_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_20_io_in_kv = local_pes_27_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_20_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_20_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_20_io_in_stage = local_pes_28_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_21_clock = clock;
  assign local_pes_28_21_reset = reset;
  assign local_pes_28_21_io_in_q = local_pes_28_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_21_io_in_sum = local_pes_28_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_21_io_in_sum_exp = local_pes_28_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_21_io_in_kv = local_pes_27_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_21_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_21_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_21_io_in_stage = local_pes_28_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_22_clock = clock;
  assign local_pes_28_22_reset = reset;
  assign local_pes_28_22_io_in_q = local_pes_28_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_22_io_in_sum = local_pes_28_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_22_io_in_sum_exp = local_pes_28_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_22_io_in_kv = local_pes_27_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_22_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_22_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_22_io_in_stage = local_pes_28_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_23_clock = clock;
  assign local_pes_28_23_reset = reset;
  assign local_pes_28_23_io_in_q = local_pes_28_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_23_io_in_sum = local_pes_28_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_23_io_in_sum_exp = local_pes_28_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_23_io_in_kv = local_pes_27_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_23_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_23_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_23_io_in_stage = local_pes_28_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_24_clock = clock;
  assign local_pes_28_24_reset = reset;
  assign local_pes_28_24_io_in_q = local_pes_28_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_24_io_in_sum = local_pes_28_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_24_io_in_sum_exp = local_pes_28_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_24_io_in_kv = local_pes_27_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_24_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_24_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_24_io_in_stage = local_pes_28_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_25_clock = clock;
  assign local_pes_28_25_reset = reset;
  assign local_pes_28_25_io_in_q = local_pes_28_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_25_io_in_sum = local_pes_28_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_25_io_in_sum_exp = local_pes_28_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_25_io_in_kv = local_pes_27_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_25_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_25_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_25_io_in_stage = local_pes_28_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_26_clock = clock;
  assign local_pes_28_26_reset = reset;
  assign local_pes_28_26_io_in_q = local_pes_28_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_26_io_in_sum = local_pes_28_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_26_io_in_sum_exp = local_pes_28_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_26_io_in_kv = local_pes_27_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_26_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_26_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_26_io_in_stage = local_pes_28_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_27_clock = clock;
  assign local_pes_28_27_reset = reset;
  assign local_pes_28_27_io_in_q = local_pes_28_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_27_io_in_sum = local_pes_28_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_27_io_in_sum_exp = local_pes_28_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_27_io_in_kv = local_pes_27_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_27_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_27_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_27_io_in_stage = local_pes_28_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_28_clock = clock;
  assign local_pes_28_28_reset = reset;
  assign local_pes_28_28_io_in_q = local_pes_28_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_28_io_in_sum = local_pes_28_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_28_io_in_sum_exp = local_pes_28_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_28_io_in_kv = local_pes_27_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_28_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_28_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_28_io_in_stage = local_pes_28_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_29_clock = clock;
  assign local_pes_28_29_reset = reset;
  assign local_pes_28_29_io_in_q = local_pes_28_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_29_io_in_sum = local_pes_28_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_29_io_in_sum_exp = local_pes_28_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_29_io_in_kv = local_pes_27_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_29_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_29_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_29_io_in_stage = local_pes_28_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_30_clock = clock;
  assign local_pes_28_30_reset = reset;
  assign local_pes_28_30_io_in_q = local_pes_28_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_30_io_in_sum = local_pes_28_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_30_io_in_sum_exp = local_pes_28_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_30_io_in_kv = local_pes_27_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_30_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_30_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_30_io_in_stage = local_pes_28_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_28_31_clock = clock;
  assign local_pes_28_31_reset = reset;
  assign local_pes_28_31_io_in_q = local_pes_28_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_28_31_io_in_sum = local_pes_28_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_28_31_io_in_sum_exp = local_pes_28_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_28_31_io_in_kv = local_pes_27_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_28_31_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_28_31_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_28_31_io_in_stage = local_pes_28_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_0_clock = clock;
  assign local_pes_29_0_reset = reset;
  assign local_pes_29_0_io_in_q = io_q_ports_29; // @[PEArray.scala 51:37]
  assign local_pes_29_0_io_in_kv = io_kv_ports_60; // @[PEArray.scala 40:34]
  assign local_pes_29_0_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_0_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_0_io_in_stage = io_stage_ports_29; // @[PEArray.scala 52:41]
  assign local_pes_29_1_clock = clock;
  assign local_pes_29_1_reset = reset;
  assign local_pes_29_1_io_in_q = local_pes_29_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_1_io_in_sum = local_pes_29_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_29_1_io_in_kv = local_pes_28_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_1_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_1_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_1_io_in_stage = local_pes_29_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_2_clock = clock;
  assign local_pes_29_2_reset = reset;
  assign local_pes_29_2_io_in_q = local_pes_29_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_2_io_in_sum = local_pes_29_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_2_io_in_sum_exp = local_pes_29_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_2_io_in_kv = local_pes_28_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_2_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_2_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_2_io_in_stage = local_pes_29_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_3_clock = clock;
  assign local_pes_29_3_reset = reset;
  assign local_pes_29_3_io_in_q = local_pes_29_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_3_io_in_sum = local_pes_29_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_3_io_in_sum_exp = local_pes_29_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_3_io_in_kv = local_pes_28_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_3_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_3_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_3_io_in_stage = local_pes_29_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_4_clock = clock;
  assign local_pes_29_4_reset = reset;
  assign local_pes_29_4_io_in_q = local_pes_29_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_4_io_in_sum = local_pes_29_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_4_io_in_sum_exp = local_pes_29_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_4_io_in_kv = local_pes_28_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_4_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_4_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_4_io_in_stage = local_pes_29_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_5_clock = clock;
  assign local_pes_29_5_reset = reset;
  assign local_pes_29_5_io_in_q = local_pes_29_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_5_io_in_sum = local_pes_29_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_5_io_in_sum_exp = local_pes_29_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_5_io_in_kv = local_pes_28_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_5_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_5_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_5_io_in_stage = local_pes_29_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_6_clock = clock;
  assign local_pes_29_6_reset = reset;
  assign local_pes_29_6_io_in_q = local_pes_29_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_6_io_in_sum = local_pes_29_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_6_io_in_sum_exp = local_pes_29_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_6_io_in_kv = local_pes_28_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_6_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_6_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_6_io_in_stage = local_pes_29_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_7_clock = clock;
  assign local_pes_29_7_reset = reset;
  assign local_pes_29_7_io_in_q = local_pes_29_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_7_io_in_sum = local_pes_29_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_7_io_in_sum_exp = local_pes_29_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_7_io_in_kv = local_pes_28_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_7_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_7_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_7_io_in_stage = local_pes_29_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_8_clock = clock;
  assign local_pes_29_8_reset = reset;
  assign local_pes_29_8_io_in_q = local_pes_29_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_8_io_in_sum = local_pes_29_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_8_io_in_sum_exp = local_pes_29_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_8_io_in_kv = local_pes_28_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_8_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_8_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_8_io_in_stage = local_pes_29_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_9_clock = clock;
  assign local_pes_29_9_reset = reset;
  assign local_pes_29_9_io_in_q = local_pes_29_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_9_io_in_sum = local_pes_29_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_9_io_in_sum_exp = local_pes_29_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_9_io_in_kv = local_pes_28_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_9_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_9_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_9_io_in_stage = local_pes_29_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_10_clock = clock;
  assign local_pes_29_10_reset = reset;
  assign local_pes_29_10_io_in_q = local_pes_29_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_10_io_in_sum = local_pes_29_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_10_io_in_sum_exp = local_pes_29_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_10_io_in_kv = local_pes_28_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_10_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_10_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_10_io_in_stage = local_pes_29_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_11_clock = clock;
  assign local_pes_29_11_reset = reset;
  assign local_pes_29_11_io_in_q = local_pes_29_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_11_io_in_sum = local_pes_29_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_11_io_in_sum_exp = local_pes_29_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_11_io_in_kv = local_pes_28_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_11_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_11_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_11_io_in_stage = local_pes_29_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_12_clock = clock;
  assign local_pes_29_12_reset = reset;
  assign local_pes_29_12_io_in_q = local_pes_29_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_12_io_in_sum = local_pes_29_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_12_io_in_sum_exp = local_pes_29_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_12_io_in_kv = local_pes_28_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_12_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_12_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_12_io_in_stage = local_pes_29_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_13_clock = clock;
  assign local_pes_29_13_reset = reset;
  assign local_pes_29_13_io_in_q = local_pes_29_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_13_io_in_sum = local_pes_29_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_13_io_in_sum_exp = local_pes_29_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_13_io_in_kv = local_pes_28_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_13_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_13_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_13_io_in_stage = local_pes_29_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_14_clock = clock;
  assign local_pes_29_14_reset = reset;
  assign local_pes_29_14_io_in_q = local_pes_29_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_14_io_in_sum = local_pes_29_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_14_io_in_sum_exp = local_pes_29_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_14_io_in_kv = local_pes_28_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_14_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_14_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_14_io_in_stage = local_pes_29_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_15_clock = clock;
  assign local_pes_29_15_reset = reset;
  assign local_pes_29_15_io_in_q = local_pes_29_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_15_io_in_sum = local_pes_29_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_15_io_in_sum_exp = local_pes_29_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_15_io_in_kv = local_pes_28_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_15_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_15_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_15_io_in_stage = local_pes_29_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_16_clock = clock;
  assign local_pes_29_16_reset = reset;
  assign local_pes_29_16_io_in_q = local_pes_29_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_16_io_in_sum = local_pes_29_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_16_io_in_sum_exp = local_pes_29_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_16_io_in_kv = local_pes_28_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_16_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_16_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_16_io_in_stage = local_pes_29_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_17_clock = clock;
  assign local_pes_29_17_reset = reset;
  assign local_pes_29_17_io_in_q = local_pes_29_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_17_io_in_sum = local_pes_29_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_17_io_in_sum_exp = local_pes_29_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_17_io_in_kv = local_pes_28_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_17_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_17_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_17_io_in_stage = local_pes_29_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_18_clock = clock;
  assign local_pes_29_18_reset = reset;
  assign local_pes_29_18_io_in_q = local_pes_29_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_18_io_in_sum = local_pes_29_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_18_io_in_sum_exp = local_pes_29_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_18_io_in_kv = local_pes_28_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_18_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_18_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_18_io_in_stage = local_pes_29_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_19_clock = clock;
  assign local_pes_29_19_reset = reset;
  assign local_pes_29_19_io_in_q = local_pes_29_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_19_io_in_sum = local_pes_29_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_19_io_in_sum_exp = local_pes_29_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_19_io_in_kv = local_pes_28_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_19_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_19_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_19_io_in_stage = local_pes_29_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_20_clock = clock;
  assign local_pes_29_20_reset = reset;
  assign local_pes_29_20_io_in_q = local_pes_29_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_20_io_in_sum = local_pes_29_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_20_io_in_sum_exp = local_pes_29_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_20_io_in_kv = local_pes_28_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_20_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_20_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_20_io_in_stage = local_pes_29_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_21_clock = clock;
  assign local_pes_29_21_reset = reset;
  assign local_pes_29_21_io_in_q = local_pes_29_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_21_io_in_sum = local_pes_29_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_21_io_in_sum_exp = local_pes_29_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_21_io_in_kv = local_pes_28_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_21_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_21_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_21_io_in_stage = local_pes_29_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_22_clock = clock;
  assign local_pes_29_22_reset = reset;
  assign local_pes_29_22_io_in_q = local_pes_29_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_22_io_in_sum = local_pes_29_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_22_io_in_sum_exp = local_pes_29_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_22_io_in_kv = local_pes_28_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_22_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_22_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_22_io_in_stage = local_pes_29_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_23_clock = clock;
  assign local_pes_29_23_reset = reset;
  assign local_pes_29_23_io_in_q = local_pes_29_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_23_io_in_sum = local_pes_29_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_23_io_in_sum_exp = local_pes_29_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_23_io_in_kv = local_pes_28_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_23_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_23_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_23_io_in_stage = local_pes_29_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_24_clock = clock;
  assign local_pes_29_24_reset = reset;
  assign local_pes_29_24_io_in_q = local_pes_29_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_24_io_in_sum = local_pes_29_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_24_io_in_sum_exp = local_pes_29_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_24_io_in_kv = local_pes_28_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_24_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_24_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_24_io_in_stage = local_pes_29_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_25_clock = clock;
  assign local_pes_29_25_reset = reset;
  assign local_pes_29_25_io_in_q = local_pes_29_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_25_io_in_sum = local_pes_29_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_25_io_in_sum_exp = local_pes_29_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_25_io_in_kv = local_pes_28_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_25_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_25_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_25_io_in_stage = local_pes_29_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_26_clock = clock;
  assign local_pes_29_26_reset = reset;
  assign local_pes_29_26_io_in_q = local_pes_29_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_26_io_in_sum = local_pes_29_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_26_io_in_sum_exp = local_pes_29_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_26_io_in_kv = local_pes_28_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_26_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_26_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_26_io_in_stage = local_pes_29_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_27_clock = clock;
  assign local_pes_29_27_reset = reset;
  assign local_pes_29_27_io_in_q = local_pes_29_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_27_io_in_sum = local_pes_29_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_27_io_in_sum_exp = local_pes_29_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_27_io_in_kv = local_pes_28_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_27_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_27_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_27_io_in_stage = local_pes_29_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_28_clock = clock;
  assign local_pes_29_28_reset = reset;
  assign local_pes_29_28_io_in_q = local_pes_29_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_28_io_in_sum = local_pes_29_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_28_io_in_sum_exp = local_pes_29_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_28_io_in_kv = local_pes_28_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_28_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_28_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_28_io_in_stage = local_pes_29_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_29_clock = clock;
  assign local_pes_29_29_reset = reset;
  assign local_pes_29_29_io_in_q = local_pes_29_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_29_io_in_sum = local_pes_29_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_29_io_in_sum_exp = local_pes_29_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_29_io_in_kv = local_pes_28_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_29_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_29_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_29_io_in_stage = local_pes_29_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_30_clock = clock;
  assign local_pes_29_30_reset = reset;
  assign local_pes_29_30_io_in_q = local_pes_29_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_30_io_in_sum = local_pes_29_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_30_io_in_sum_exp = local_pes_29_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_30_io_in_kv = local_pes_28_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_30_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_30_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_30_io_in_stage = local_pes_29_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_29_31_clock = clock;
  assign local_pes_29_31_reset = reset;
  assign local_pes_29_31_io_in_q = local_pes_29_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_29_31_io_in_sum = local_pes_29_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_29_31_io_in_sum_exp = local_pes_29_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_29_31_io_in_kv = local_pes_28_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_29_31_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_29_31_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_29_31_io_in_stage = local_pes_29_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_0_clock = clock;
  assign local_pes_30_0_reset = reset;
  assign local_pes_30_0_io_in_q = io_q_ports_30; // @[PEArray.scala 51:37]
  assign local_pes_30_0_io_in_kv = io_kv_ports_61; // @[PEArray.scala 40:34]
  assign local_pes_30_0_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_0_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_0_io_in_stage = io_stage_ports_30; // @[PEArray.scala 52:41]
  assign local_pes_30_1_clock = clock;
  assign local_pes_30_1_reset = reset;
  assign local_pes_30_1_io_in_q = local_pes_30_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_1_io_in_sum = local_pes_30_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_30_1_io_in_kv = local_pes_29_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_1_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_1_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_1_io_in_stage = local_pes_30_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_2_clock = clock;
  assign local_pes_30_2_reset = reset;
  assign local_pes_30_2_io_in_q = local_pes_30_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_2_io_in_sum = local_pes_30_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_2_io_in_sum_exp = local_pes_30_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_2_io_in_kv = local_pes_29_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_2_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_2_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_2_io_in_stage = local_pes_30_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_3_clock = clock;
  assign local_pes_30_3_reset = reset;
  assign local_pes_30_3_io_in_q = local_pes_30_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_3_io_in_sum = local_pes_30_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_3_io_in_sum_exp = local_pes_30_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_3_io_in_kv = local_pes_29_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_3_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_3_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_3_io_in_stage = local_pes_30_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_4_clock = clock;
  assign local_pes_30_4_reset = reset;
  assign local_pes_30_4_io_in_q = local_pes_30_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_4_io_in_sum = local_pes_30_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_4_io_in_sum_exp = local_pes_30_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_4_io_in_kv = local_pes_29_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_4_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_4_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_4_io_in_stage = local_pes_30_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_5_clock = clock;
  assign local_pes_30_5_reset = reset;
  assign local_pes_30_5_io_in_q = local_pes_30_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_5_io_in_sum = local_pes_30_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_5_io_in_sum_exp = local_pes_30_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_5_io_in_kv = local_pes_29_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_5_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_5_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_5_io_in_stage = local_pes_30_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_6_clock = clock;
  assign local_pes_30_6_reset = reset;
  assign local_pes_30_6_io_in_q = local_pes_30_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_6_io_in_sum = local_pes_30_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_6_io_in_sum_exp = local_pes_30_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_6_io_in_kv = local_pes_29_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_6_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_6_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_6_io_in_stage = local_pes_30_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_7_clock = clock;
  assign local_pes_30_7_reset = reset;
  assign local_pes_30_7_io_in_q = local_pes_30_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_7_io_in_sum = local_pes_30_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_7_io_in_sum_exp = local_pes_30_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_7_io_in_kv = local_pes_29_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_7_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_7_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_7_io_in_stage = local_pes_30_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_8_clock = clock;
  assign local_pes_30_8_reset = reset;
  assign local_pes_30_8_io_in_q = local_pes_30_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_8_io_in_sum = local_pes_30_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_8_io_in_sum_exp = local_pes_30_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_8_io_in_kv = local_pes_29_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_8_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_8_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_8_io_in_stage = local_pes_30_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_9_clock = clock;
  assign local_pes_30_9_reset = reset;
  assign local_pes_30_9_io_in_q = local_pes_30_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_9_io_in_sum = local_pes_30_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_9_io_in_sum_exp = local_pes_30_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_9_io_in_kv = local_pes_29_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_9_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_9_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_9_io_in_stage = local_pes_30_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_10_clock = clock;
  assign local_pes_30_10_reset = reset;
  assign local_pes_30_10_io_in_q = local_pes_30_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_10_io_in_sum = local_pes_30_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_10_io_in_sum_exp = local_pes_30_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_10_io_in_kv = local_pes_29_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_10_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_10_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_10_io_in_stage = local_pes_30_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_11_clock = clock;
  assign local_pes_30_11_reset = reset;
  assign local_pes_30_11_io_in_q = local_pes_30_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_11_io_in_sum = local_pes_30_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_11_io_in_sum_exp = local_pes_30_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_11_io_in_kv = local_pes_29_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_11_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_11_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_11_io_in_stage = local_pes_30_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_12_clock = clock;
  assign local_pes_30_12_reset = reset;
  assign local_pes_30_12_io_in_q = local_pes_30_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_12_io_in_sum = local_pes_30_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_12_io_in_sum_exp = local_pes_30_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_12_io_in_kv = local_pes_29_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_12_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_12_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_12_io_in_stage = local_pes_30_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_13_clock = clock;
  assign local_pes_30_13_reset = reset;
  assign local_pes_30_13_io_in_q = local_pes_30_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_13_io_in_sum = local_pes_30_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_13_io_in_sum_exp = local_pes_30_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_13_io_in_kv = local_pes_29_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_13_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_13_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_13_io_in_stage = local_pes_30_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_14_clock = clock;
  assign local_pes_30_14_reset = reset;
  assign local_pes_30_14_io_in_q = local_pes_30_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_14_io_in_sum = local_pes_30_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_14_io_in_sum_exp = local_pes_30_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_14_io_in_kv = local_pes_29_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_14_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_14_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_14_io_in_stage = local_pes_30_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_15_clock = clock;
  assign local_pes_30_15_reset = reset;
  assign local_pes_30_15_io_in_q = local_pes_30_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_15_io_in_sum = local_pes_30_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_15_io_in_sum_exp = local_pes_30_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_15_io_in_kv = local_pes_29_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_15_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_15_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_15_io_in_stage = local_pes_30_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_16_clock = clock;
  assign local_pes_30_16_reset = reset;
  assign local_pes_30_16_io_in_q = local_pes_30_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_16_io_in_sum = local_pes_30_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_16_io_in_sum_exp = local_pes_30_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_16_io_in_kv = local_pes_29_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_16_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_16_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_16_io_in_stage = local_pes_30_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_17_clock = clock;
  assign local_pes_30_17_reset = reset;
  assign local_pes_30_17_io_in_q = local_pes_30_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_17_io_in_sum = local_pes_30_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_17_io_in_sum_exp = local_pes_30_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_17_io_in_kv = local_pes_29_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_17_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_17_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_17_io_in_stage = local_pes_30_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_18_clock = clock;
  assign local_pes_30_18_reset = reset;
  assign local_pes_30_18_io_in_q = local_pes_30_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_18_io_in_sum = local_pes_30_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_18_io_in_sum_exp = local_pes_30_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_18_io_in_kv = local_pes_29_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_18_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_18_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_18_io_in_stage = local_pes_30_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_19_clock = clock;
  assign local_pes_30_19_reset = reset;
  assign local_pes_30_19_io_in_q = local_pes_30_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_19_io_in_sum = local_pes_30_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_19_io_in_sum_exp = local_pes_30_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_19_io_in_kv = local_pes_29_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_19_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_19_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_19_io_in_stage = local_pes_30_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_20_clock = clock;
  assign local_pes_30_20_reset = reset;
  assign local_pes_30_20_io_in_q = local_pes_30_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_20_io_in_sum = local_pes_30_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_20_io_in_sum_exp = local_pes_30_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_20_io_in_kv = local_pes_29_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_20_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_20_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_20_io_in_stage = local_pes_30_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_21_clock = clock;
  assign local_pes_30_21_reset = reset;
  assign local_pes_30_21_io_in_q = local_pes_30_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_21_io_in_sum = local_pes_30_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_21_io_in_sum_exp = local_pes_30_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_21_io_in_kv = local_pes_29_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_21_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_21_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_21_io_in_stage = local_pes_30_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_22_clock = clock;
  assign local_pes_30_22_reset = reset;
  assign local_pes_30_22_io_in_q = local_pes_30_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_22_io_in_sum = local_pes_30_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_22_io_in_sum_exp = local_pes_30_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_22_io_in_kv = local_pes_29_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_22_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_22_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_22_io_in_stage = local_pes_30_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_23_clock = clock;
  assign local_pes_30_23_reset = reset;
  assign local_pes_30_23_io_in_q = local_pes_30_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_23_io_in_sum = local_pes_30_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_23_io_in_sum_exp = local_pes_30_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_23_io_in_kv = local_pes_29_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_23_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_23_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_23_io_in_stage = local_pes_30_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_24_clock = clock;
  assign local_pes_30_24_reset = reset;
  assign local_pes_30_24_io_in_q = local_pes_30_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_24_io_in_sum = local_pes_30_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_24_io_in_sum_exp = local_pes_30_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_24_io_in_kv = local_pes_29_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_24_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_24_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_24_io_in_stage = local_pes_30_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_25_clock = clock;
  assign local_pes_30_25_reset = reset;
  assign local_pes_30_25_io_in_q = local_pes_30_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_25_io_in_sum = local_pes_30_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_25_io_in_sum_exp = local_pes_30_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_25_io_in_kv = local_pes_29_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_25_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_25_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_25_io_in_stage = local_pes_30_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_26_clock = clock;
  assign local_pes_30_26_reset = reset;
  assign local_pes_30_26_io_in_q = local_pes_30_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_26_io_in_sum = local_pes_30_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_26_io_in_sum_exp = local_pes_30_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_26_io_in_kv = local_pes_29_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_26_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_26_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_26_io_in_stage = local_pes_30_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_27_clock = clock;
  assign local_pes_30_27_reset = reset;
  assign local_pes_30_27_io_in_q = local_pes_30_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_27_io_in_sum = local_pes_30_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_27_io_in_sum_exp = local_pes_30_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_27_io_in_kv = local_pes_29_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_27_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_27_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_27_io_in_stage = local_pes_30_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_28_clock = clock;
  assign local_pes_30_28_reset = reset;
  assign local_pes_30_28_io_in_q = local_pes_30_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_28_io_in_sum = local_pes_30_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_28_io_in_sum_exp = local_pes_30_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_28_io_in_kv = local_pes_29_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_28_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_28_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_28_io_in_stage = local_pes_30_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_29_clock = clock;
  assign local_pes_30_29_reset = reset;
  assign local_pes_30_29_io_in_q = local_pes_30_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_29_io_in_sum = local_pes_30_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_29_io_in_sum_exp = local_pes_30_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_29_io_in_kv = local_pes_29_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_29_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_29_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_29_io_in_stage = local_pes_30_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_30_clock = clock;
  assign local_pes_30_30_reset = reset;
  assign local_pes_30_30_io_in_q = local_pes_30_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_30_io_in_sum = local_pes_30_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_30_io_in_sum_exp = local_pes_30_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_30_io_in_kv = local_pes_29_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_30_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_30_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_30_io_in_stage = local_pes_30_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_30_31_clock = clock;
  assign local_pes_30_31_reset = reset;
  assign local_pes_30_31_io_in_q = local_pes_30_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_30_31_io_in_sum = local_pes_30_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_30_31_io_in_sum_exp = local_pes_30_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_30_31_io_in_kv = local_pes_29_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_30_31_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_30_31_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_30_31_io_in_stage = local_pes_30_30_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_0_clock = clock;
  assign local_pes_31_0_reset = reset;
  assign local_pes_31_0_io_in_q = io_q_ports_31; // @[PEArray.scala 51:37]
  assign local_pes_31_0_io_in_kv = io_kv_ports_62; // @[PEArray.scala 40:34]
  assign local_pes_31_0_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_0_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_0_io_in_stage = io_stage_ports_31; // @[PEArray.scala 52:41]
  assign local_pes_31_1_clock = clock;
  assign local_pes_31_1_reset = reset;
  assign local_pes_31_1_io_in_q = local_pes_31_0_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_1_io_in_sum = local_pes_31_0_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 54:43]
  assign local_pes_31_1_io_in_kv = local_pes_30_0_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_1_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_1_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_1_io_in_stage = local_pes_31_0_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_2_clock = clock;
  assign local_pes_31_2_reset = reset;
  assign local_pes_31_2_io_in_q = local_pes_31_1_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_2_io_in_sum = local_pes_31_1_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_2_io_in_sum_exp = local_pes_31_1_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_2_io_in_kv = local_pes_30_1_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_2_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_2_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_2_io_in_stage = local_pes_31_1_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_3_clock = clock;
  assign local_pes_31_3_reset = reset;
  assign local_pes_31_3_io_in_q = local_pes_31_2_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_3_io_in_sum = local_pes_31_2_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_3_io_in_sum_exp = local_pes_31_2_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_3_io_in_kv = local_pes_30_2_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_3_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_3_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_3_io_in_stage = local_pes_31_2_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_4_clock = clock;
  assign local_pes_31_4_reset = reset;
  assign local_pes_31_4_io_in_q = local_pes_31_3_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_4_io_in_sum = local_pes_31_3_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_4_io_in_sum_exp = local_pes_31_3_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_4_io_in_kv = local_pes_30_3_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_4_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_4_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_4_io_in_stage = local_pes_31_3_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_5_clock = clock;
  assign local_pes_31_5_reset = reset;
  assign local_pes_31_5_io_in_q = local_pes_31_4_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_5_io_in_sum = local_pes_31_4_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_5_io_in_sum_exp = local_pes_31_4_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_5_io_in_kv = local_pes_30_4_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_5_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_5_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_5_io_in_stage = local_pes_31_4_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_6_clock = clock;
  assign local_pes_31_6_reset = reset;
  assign local_pes_31_6_io_in_q = local_pes_31_5_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_6_io_in_sum = local_pes_31_5_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_6_io_in_sum_exp = local_pes_31_5_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_6_io_in_kv = local_pes_30_5_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_6_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_6_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_6_io_in_stage = local_pes_31_5_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_7_clock = clock;
  assign local_pes_31_7_reset = reset;
  assign local_pes_31_7_io_in_q = local_pes_31_6_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_7_io_in_sum = local_pes_31_6_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_7_io_in_sum_exp = local_pes_31_6_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_7_io_in_kv = local_pes_30_6_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_7_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_7_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_7_io_in_stage = local_pes_31_6_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_8_clock = clock;
  assign local_pes_31_8_reset = reset;
  assign local_pes_31_8_io_in_q = local_pes_31_7_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_8_io_in_sum = local_pes_31_7_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_8_io_in_sum_exp = local_pes_31_7_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_8_io_in_kv = local_pes_30_7_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_8_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_8_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_8_io_in_stage = local_pes_31_7_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_9_clock = clock;
  assign local_pes_31_9_reset = reset;
  assign local_pes_31_9_io_in_q = local_pes_31_8_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_9_io_in_sum = local_pes_31_8_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_9_io_in_sum_exp = local_pes_31_8_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_9_io_in_kv = local_pes_30_8_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_9_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_9_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_9_io_in_stage = local_pes_31_8_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_10_clock = clock;
  assign local_pes_31_10_reset = reset;
  assign local_pes_31_10_io_in_q = local_pes_31_9_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_10_io_in_sum = local_pes_31_9_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_10_io_in_sum_exp = local_pes_31_9_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_10_io_in_kv = local_pes_30_9_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_10_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_10_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_10_io_in_stage = local_pes_31_9_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_11_clock = clock;
  assign local_pes_31_11_reset = reset;
  assign local_pes_31_11_io_in_q = local_pes_31_10_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_11_io_in_sum = local_pes_31_10_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_11_io_in_sum_exp = local_pes_31_10_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_11_io_in_kv = local_pes_30_10_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_11_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_11_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_11_io_in_stage = local_pes_31_10_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_12_clock = clock;
  assign local_pes_31_12_reset = reset;
  assign local_pes_31_12_io_in_q = local_pes_31_11_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_12_io_in_sum = local_pes_31_11_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_12_io_in_sum_exp = local_pes_31_11_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_12_io_in_kv = local_pes_30_11_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_12_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_12_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_12_io_in_stage = local_pes_31_11_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_13_clock = clock;
  assign local_pes_31_13_reset = reset;
  assign local_pes_31_13_io_in_q = local_pes_31_12_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_13_io_in_sum = local_pes_31_12_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_13_io_in_sum_exp = local_pes_31_12_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_13_io_in_kv = local_pes_30_12_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_13_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_13_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_13_io_in_stage = local_pes_31_12_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_14_clock = clock;
  assign local_pes_31_14_reset = reset;
  assign local_pes_31_14_io_in_q = local_pes_31_13_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_14_io_in_sum = local_pes_31_13_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_14_io_in_sum_exp = local_pes_31_13_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_14_io_in_kv = local_pes_30_13_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_14_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_14_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_14_io_in_stage = local_pes_31_13_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_15_clock = clock;
  assign local_pes_31_15_reset = reset;
  assign local_pes_31_15_io_in_q = local_pes_31_14_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_15_io_in_sum = local_pes_31_14_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_15_io_in_sum_exp = local_pes_31_14_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_15_io_in_kv = local_pes_30_14_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_15_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_15_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_15_io_in_stage = local_pes_31_14_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_16_clock = clock;
  assign local_pes_31_16_reset = reset;
  assign local_pes_31_16_io_in_q = local_pes_31_15_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_16_io_in_sum = local_pes_31_15_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_16_io_in_sum_exp = local_pes_31_15_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_16_io_in_kv = local_pes_30_15_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_16_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_16_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_16_io_in_stage = local_pes_31_15_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_17_clock = clock;
  assign local_pes_31_17_reset = reset;
  assign local_pes_31_17_io_in_q = local_pes_31_16_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_17_io_in_sum = local_pes_31_16_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_17_io_in_sum_exp = local_pes_31_16_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_17_io_in_kv = local_pes_30_16_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_17_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_17_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_17_io_in_stage = local_pes_31_16_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_18_clock = clock;
  assign local_pes_31_18_reset = reset;
  assign local_pes_31_18_io_in_q = local_pes_31_17_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_18_io_in_sum = local_pes_31_17_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_18_io_in_sum_exp = local_pes_31_17_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_18_io_in_kv = local_pes_30_17_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_18_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_18_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_18_io_in_stage = local_pes_31_17_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_19_clock = clock;
  assign local_pes_31_19_reset = reset;
  assign local_pes_31_19_io_in_q = local_pes_31_18_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_19_io_in_sum = local_pes_31_18_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_19_io_in_sum_exp = local_pes_31_18_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_19_io_in_kv = local_pes_30_18_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_19_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_19_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_19_io_in_stage = local_pes_31_18_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_20_clock = clock;
  assign local_pes_31_20_reset = reset;
  assign local_pes_31_20_io_in_q = local_pes_31_19_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_20_io_in_sum = local_pes_31_19_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_20_io_in_sum_exp = local_pes_31_19_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_20_io_in_kv = local_pes_30_19_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_20_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_20_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_20_io_in_stage = local_pes_31_19_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_21_clock = clock;
  assign local_pes_31_21_reset = reset;
  assign local_pes_31_21_io_in_q = local_pes_31_20_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_21_io_in_sum = local_pes_31_20_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_21_io_in_sum_exp = local_pes_31_20_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_21_io_in_kv = local_pes_30_20_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_21_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_21_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_21_io_in_stage = local_pes_31_20_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_22_clock = clock;
  assign local_pes_31_22_reset = reset;
  assign local_pes_31_22_io_in_q = local_pes_31_21_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_22_io_in_sum = local_pes_31_21_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_22_io_in_sum_exp = local_pes_31_21_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_22_io_in_kv = local_pes_30_21_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_22_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_22_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_22_io_in_stage = local_pes_31_21_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_23_clock = clock;
  assign local_pes_31_23_reset = reset;
  assign local_pes_31_23_io_in_q = local_pes_31_22_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_23_io_in_sum = local_pes_31_22_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_23_io_in_sum_exp = local_pes_31_22_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_23_io_in_kv = local_pes_30_22_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_23_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_23_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_23_io_in_stage = local_pes_31_22_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_24_clock = clock;
  assign local_pes_31_24_reset = reset;
  assign local_pes_31_24_io_in_q = local_pes_31_23_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_24_io_in_sum = local_pes_31_23_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_24_io_in_sum_exp = local_pes_31_23_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_24_io_in_kv = local_pes_30_23_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_24_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_24_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_24_io_in_stage = local_pes_31_23_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_25_clock = clock;
  assign local_pes_31_25_reset = reset;
  assign local_pes_31_25_io_in_q = local_pes_31_24_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_25_io_in_sum = local_pes_31_24_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_25_io_in_sum_exp = local_pes_31_24_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_25_io_in_kv = local_pes_30_24_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_25_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_25_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_25_io_in_stage = local_pes_31_24_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_26_clock = clock;
  assign local_pes_31_26_reset = reset;
  assign local_pes_31_26_io_in_q = local_pes_31_25_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_26_io_in_sum = local_pes_31_25_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_26_io_in_sum_exp = local_pes_31_25_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_26_io_in_kv = local_pes_30_25_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_26_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_26_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_26_io_in_stage = local_pes_31_25_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_27_clock = clock;
  assign local_pes_31_27_reset = reset;
  assign local_pes_31_27_io_in_q = local_pes_31_26_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_27_io_in_sum = local_pes_31_26_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_27_io_in_sum_exp = local_pes_31_26_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_27_io_in_kv = local_pes_30_26_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_27_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_27_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_27_io_in_stage = local_pes_31_26_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_28_clock = clock;
  assign local_pes_31_28_reset = reset;
  assign local_pes_31_28_io_in_q = local_pes_31_27_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_28_io_in_sum = local_pes_31_27_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_28_io_in_sum_exp = local_pes_31_27_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_28_io_in_kv = local_pes_30_27_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_28_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_28_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_28_io_in_stage = local_pes_31_27_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_29_clock = clock;
  assign local_pes_31_29_reset = reset;
  assign local_pes_31_29_io_in_q = local_pes_31_28_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_29_io_in_sum = local_pes_31_28_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_29_io_in_sum_exp = local_pes_31_28_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_29_io_in_kv = local_pes_30_28_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_29_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_29_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_29_io_in_stage = local_pes_31_28_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_30_clock = clock;
  assign local_pes_31_30_reset = reset;
  assign local_pes_31_30_io_in_q = local_pes_31_29_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_30_io_in_sum = local_pes_31_29_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_30_io_in_sum_exp = local_pes_31_29_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_30_io_in_kv = local_pes_30_29_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_30_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_30_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_30_io_in_stage = local_pes_31_29_io_out_stage; // @[PEArray.scala 52:41]
  assign local_pes_31_31_clock = clock;
  assign local_pes_31_31_reset = reset;
  assign local_pes_31_31_io_in_q = local_pes_31_30_io_out_q; // @[PEArray.scala 51:37]
  assign local_pes_31_31_io_in_sum = local_pes_31_30_io_out_sum; // @[PEArray.scala 53:39]
  assign local_pes_31_31_io_in_sum_exp = local_pes_31_30_io_out_sum_exp; // @[PEArray.scala 54:43]
  assign local_pes_31_31_io_in_kv = local_pes_30_30_io_out_kv; // @[PEArray.scala 45:38]
  assign local_pes_31_31_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 56:47]
  assign local_pes_31_31_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 55:43]
  assign local_pes_31_31_io_in_stage = local_pes_31_30_io_out_stage; // @[PEArray.scala 52:41]
  assign global_col_pes_0_0_clock = clock;
  assign global_col_pes_0_0_reset = reset;
  assign global_col_pes_0_0_io_in_q = local_pes_0_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_0_0_io_in_sum = local_pes_0_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_0_0_io_in_sum_exp = local_pes_0_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_0_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_0_0_io_in_inv_sum_exp = inv_modules_0_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_0_0_io_in_inv_sum = _GEN_0[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_0_0_io_in_stage = local_pes_0_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_1_0_clock = clock;
  assign global_col_pes_1_0_reset = reset;
  assign global_col_pes_1_0_io_in_q = local_pes_1_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_1_0_io_in_sum = local_pes_1_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_1_0_io_in_sum_exp = local_pes_1_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_1_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_1_0_io_in_inv_sum_exp = inv_modules_1_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_1_0_io_in_inv_sum = _GEN_64[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_1_0_io_in_stage = local_pes_1_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_2_0_clock = clock;
  assign global_col_pes_2_0_reset = reset;
  assign global_col_pes_2_0_io_in_q = local_pes_2_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_2_0_io_in_sum = local_pes_2_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_2_0_io_in_sum_exp = local_pes_2_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_2_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_2_0_io_in_inv_sum_exp = inv_modules_2_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_2_0_io_in_inv_sum = _GEN_128[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_2_0_io_in_stage = local_pes_2_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_3_0_clock = clock;
  assign global_col_pes_3_0_reset = reset;
  assign global_col_pes_3_0_io_in_q = local_pes_3_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_3_0_io_in_sum = local_pes_3_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_3_0_io_in_sum_exp = local_pes_3_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_3_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_3_0_io_in_inv_sum_exp = inv_modules_3_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_3_0_io_in_inv_sum = _GEN_192[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_3_0_io_in_stage = local_pes_3_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_4_0_clock = clock;
  assign global_col_pes_4_0_reset = reset;
  assign global_col_pes_4_0_io_in_q = local_pes_4_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_4_0_io_in_sum = local_pes_4_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_4_0_io_in_sum_exp = local_pes_4_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_4_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_4_0_io_in_inv_sum_exp = inv_modules_4_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_4_0_io_in_inv_sum = _GEN_256[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_4_0_io_in_stage = local_pes_4_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_5_0_clock = clock;
  assign global_col_pes_5_0_reset = reset;
  assign global_col_pes_5_0_io_in_q = local_pes_5_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_5_0_io_in_sum = local_pes_5_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_5_0_io_in_sum_exp = local_pes_5_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_5_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_5_0_io_in_inv_sum_exp = inv_modules_5_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_5_0_io_in_inv_sum = _GEN_320[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_5_0_io_in_stage = local_pes_5_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_6_0_clock = clock;
  assign global_col_pes_6_0_reset = reset;
  assign global_col_pes_6_0_io_in_q = local_pes_6_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_6_0_io_in_sum = local_pes_6_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_6_0_io_in_sum_exp = local_pes_6_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_6_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_6_0_io_in_inv_sum_exp = inv_modules_6_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_6_0_io_in_inv_sum = _GEN_384[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_6_0_io_in_stage = local_pes_6_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_7_0_clock = clock;
  assign global_col_pes_7_0_reset = reset;
  assign global_col_pes_7_0_io_in_q = local_pes_7_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_7_0_io_in_sum = local_pes_7_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_7_0_io_in_sum_exp = local_pes_7_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_7_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_7_0_io_in_inv_sum_exp = inv_modules_7_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_7_0_io_in_inv_sum = _GEN_448[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_7_0_io_in_stage = local_pes_7_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_8_0_clock = clock;
  assign global_col_pes_8_0_reset = reset;
  assign global_col_pes_8_0_io_in_q = local_pes_8_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_8_0_io_in_sum = local_pes_8_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_8_0_io_in_sum_exp = local_pes_8_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_8_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_8_0_io_in_inv_sum_exp = inv_modules_8_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_8_0_io_in_inv_sum = _GEN_512[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_8_0_io_in_stage = local_pes_8_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_9_0_clock = clock;
  assign global_col_pes_9_0_reset = reset;
  assign global_col_pes_9_0_io_in_q = local_pes_9_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_9_0_io_in_sum = local_pes_9_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_9_0_io_in_sum_exp = local_pes_9_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_9_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_9_0_io_in_inv_sum_exp = inv_modules_9_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_9_0_io_in_inv_sum = _GEN_576[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_9_0_io_in_stage = local_pes_9_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_10_0_clock = clock;
  assign global_col_pes_10_0_reset = reset;
  assign global_col_pes_10_0_io_in_q = local_pes_10_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_10_0_io_in_sum = local_pes_10_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_10_0_io_in_sum_exp = local_pes_10_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_10_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_10_0_io_in_inv_sum_exp = inv_modules_10_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_10_0_io_in_inv_sum = _GEN_640[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_10_0_io_in_stage = local_pes_10_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_11_0_clock = clock;
  assign global_col_pes_11_0_reset = reset;
  assign global_col_pes_11_0_io_in_q = local_pes_11_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_11_0_io_in_sum = local_pes_11_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_11_0_io_in_sum_exp = local_pes_11_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_11_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_11_0_io_in_inv_sum_exp = inv_modules_11_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_11_0_io_in_inv_sum = _GEN_704[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_11_0_io_in_stage = local_pes_11_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_12_0_clock = clock;
  assign global_col_pes_12_0_reset = reset;
  assign global_col_pes_12_0_io_in_q = local_pes_12_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_12_0_io_in_sum = local_pes_12_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_12_0_io_in_sum_exp = local_pes_12_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_12_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_12_0_io_in_inv_sum_exp = inv_modules_12_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_12_0_io_in_inv_sum = _GEN_768[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_12_0_io_in_stage = local_pes_12_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_13_0_clock = clock;
  assign global_col_pes_13_0_reset = reset;
  assign global_col_pes_13_0_io_in_q = local_pes_13_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_13_0_io_in_sum = local_pes_13_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_13_0_io_in_sum_exp = local_pes_13_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_13_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_13_0_io_in_inv_sum_exp = inv_modules_13_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_13_0_io_in_inv_sum = _GEN_832[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_13_0_io_in_stage = local_pes_13_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_14_0_clock = clock;
  assign global_col_pes_14_0_reset = reset;
  assign global_col_pes_14_0_io_in_q = local_pes_14_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_14_0_io_in_sum = local_pes_14_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_14_0_io_in_sum_exp = local_pes_14_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_14_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_14_0_io_in_inv_sum_exp = inv_modules_14_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_14_0_io_in_inv_sum = _GEN_896[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_14_0_io_in_stage = local_pes_14_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_15_0_clock = clock;
  assign global_col_pes_15_0_reset = reset;
  assign global_col_pes_15_0_io_in_q = local_pes_15_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_15_0_io_in_sum = local_pes_15_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_15_0_io_in_sum_exp = local_pes_15_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_15_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_15_0_io_in_inv_sum_exp = inv_modules_15_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_15_0_io_in_inv_sum = _GEN_960[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_15_0_io_in_stage = local_pes_15_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_16_0_clock = clock;
  assign global_col_pes_16_0_reset = reset;
  assign global_col_pes_16_0_io_in_q = local_pes_16_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_16_0_io_in_sum = local_pes_16_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_16_0_io_in_sum_exp = local_pes_16_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_16_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_16_0_io_in_inv_sum_exp = inv_modules_16_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_16_0_io_in_inv_sum = _GEN_1024[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_16_0_io_in_stage = local_pes_16_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_17_0_clock = clock;
  assign global_col_pes_17_0_reset = reset;
  assign global_col_pes_17_0_io_in_q = local_pes_17_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_17_0_io_in_sum = local_pes_17_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_17_0_io_in_sum_exp = local_pes_17_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_17_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_17_0_io_in_inv_sum_exp = inv_modules_17_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_17_0_io_in_inv_sum = _GEN_1088[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_17_0_io_in_stage = local_pes_17_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_18_0_clock = clock;
  assign global_col_pes_18_0_reset = reset;
  assign global_col_pes_18_0_io_in_q = local_pes_18_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_18_0_io_in_sum = local_pes_18_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_18_0_io_in_sum_exp = local_pes_18_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_18_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_18_0_io_in_inv_sum_exp = inv_modules_18_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_18_0_io_in_inv_sum = _GEN_1152[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_18_0_io_in_stage = local_pes_18_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_19_0_clock = clock;
  assign global_col_pes_19_0_reset = reset;
  assign global_col_pes_19_0_io_in_q = local_pes_19_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_19_0_io_in_sum = local_pes_19_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_19_0_io_in_sum_exp = local_pes_19_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_19_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_19_0_io_in_inv_sum_exp = inv_modules_19_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_19_0_io_in_inv_sum = _GEN_1216[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_19_0_io_in_stage = local_pes_19_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_20_0_clock = clock;
  assign global_col_pes_20_0_reset = reset;
  assign global_col_pes_20_0_io_in_q = local_pes_20_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_20_0_io_in_sum = local_pes_20_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_20_0_io_in_sum_exp = local_pes_20_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_20_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_20_0_io_in_inv_sum_exp = inv_modules_20_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_20_0_io_in_inv_sum = _GEN_1280[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_20_0_io_in_stage = local_pes_20_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_21_0_clock = clock;
  assign global_col_pes_21_0_reset = reset;
  assign global_col_pes_21_0_io_in_q = local_pes_21_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_21_0_io_in_sum = local_pes_21_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_21_0_io_in_sum_exp = local_pes_21_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_21_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_21_0_io_in_inv_sum_exp = inv_modules_21_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_21_0_io_in_inv_sum = _GEN_1344[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_21_0_io_in_stage = local_pes_21_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_22_0_clock = clock;
  assign global_col_pes_22_0_reset = reset;
  assign global_col_pes_22_0_io_in_q = local_pes_22_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_22_0_io_in_sum = local_pes_22_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_22_0_io_in_sum_exp = local_pes_22_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_22_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_22_0_io_in_inv_sum_exp = inv_modules_22_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_22_0_io_in_inv_sum = _GEN_1408[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_22_0_io_in_stage = local_pes_22_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_23_0_clock = clock;
  assign global_col_pes_23_0_reset = reset;
  assign global_col_pes_23_0_io_in_q = local_pes_23_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_23_0_io_in_sum = local_pes_23_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_23_0_io_in_sum_exp = local_pes_23_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_23_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_23_0_io_in_inv_sum_exp = inv_modules_23_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_23_0_io_in_inv_sum = _GEN_1472[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_23_0_io_in_stage = local_pes_23_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_24_0_clock = clock;
  assign global_col_pes_24_0_reset = reset;
  assign global_col_pes_24_0_io_in_q = local_pes_24_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_24_0_io_in_sum = local_pes_24_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_24_0_io_in_sum_exp = local_pes_24_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_24_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_24_0_io_in_inv_sum_exp = inv_modules_24_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_24_0_io_in_inv_sum = _GEN_1536[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_24_0_io_in_stage = local_pes_24_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_25_0_clock = clock;
  assign global_col_pes_25_0_reset = reset;
  assign global_col_pes_25_0_io_in_q = local_pes_25_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_25_0_io_in_sum = local_pes_25_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_25_0_io_in_sum_exp = local_pes_25_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_25_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_25_0_io_in_inv_sum_exp = inv_modules_25_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_25_0_io_in_inv_sum = _GEN_1600[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_25_0_io_in_stage = local_pes_25_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_26_0_clock = clock;
  assign global_col_pes_26_0_reset = reset;
  assign global_col_pes_26_0_io_in_q = local_pes_26_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_26_0_io_in_sum = local_pes_26_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_26_0_io_in_sum_exp = local_pes_26_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_26_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_26_0_io_in_inv_sum_exp = inv_modules_26_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_26_0_io_in_inv_sum = _GEN_1664[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_26_0_io_in_stage = local_pes_26_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_27_0_clock = clock;
  assign global_col_pes_27_0_reset = reset;
  assign global_col_pes_27_0_io_in_q = local_pes_27_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_27_0_io_in_sum = local_pes_27_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_27_0_io_in_sum_exp = local_pes_27_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_27_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_27_0_io_in_inv_sum_exp = inv_modules_27_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_27_0_io_in_inv_sum = _GEN_1728[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_27_0_io_in_stage = local_pes_27_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_28_0_clock = clock;
  assign global_col_pes_28_0_reset = reset;
  assign global_col_pes_28_0_io_in_q = local_pes_28_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_28_0_io_in_sum = local_pes_28_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_28_0_io_in_sum_exp = local_pes_28_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_28_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_28_0_io_in_inv_sum_exp = inv_modules_28_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_28_0_io_in_inv_sum = _GEN_1792[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_28_0_io_in_stage = local_pes_28_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_29_0_clock = clock;
  assign global_col_pes_29_0_reset = reset;
  assign global_col_pes_29_0_io_in_q = local_pes_29_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_29_0_io_in_sum = local_pes_29_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_29_0_io_in_sum_exp = local_pes_29_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_29_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_29_0_io_in_inv_sum_exp = inv_modules_29_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_29_0_io_in_inv_sum = _GEN_1856[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_29_0_io_in_stage = local_pes_29_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_30_0_clock = clock;
  assign global_col_pes_30_0_reset = reset;
  assign global_col_pes_30_0_io_in_q = local_pes_30_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_30_0_io_in_sum = local_pes_30_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_30_0_io_in_sum_exp = local_pes_30_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_30_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_30_0_io_in_inv_sum_exp = inv_modules_30_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_30_0_io_in_inv_sum = _GEN_1920[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_30_0_io_in_stage = local_pes_30_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_col_pes_31_0_clock = clock;
  assign global_col_pes_31_0_reset = reset;
  assign global_col_pes_31_0_io_in_q = local_pes_31_31_io_out_q; // @[PEArray.scala 62:42]
  assign global_col_pes_31_0_io_in_sum = local_pes_31_31_io_out_sum; // @[PEArray.scala 64:44]
  assign global_col_pes_31_0_io_in_sum_exp = local_pes_31_31_io_out_sum_exp; // @[PEArray.scala 65:48]
  assign global_col_pes_31_0_io_in_kv = io_kv_ports_63; // @[PEArray.scala 66:43]
  assign global_col_pes_31_0_io_in_inv_sum_exp = inv_modules_31_io_out_inv_sum_exp; // @[PEArray.scala 68:52]
  assign global_col_pes_31_0_io_in_inv_sum = _GEN_1984[8:0]; // @[PEArray.scala 67:48]
  assign global_col_pes_31_0_io_in_stage = local_pes_31_31_io_out_stage; // @[PEArray.scala 63:46]
  assign global_row_pes_0_0_clock = clock;
  assign global_row_pes_0_0_reset = reset;
  assign global_row_pes_0_0_io_in_q = io_q_ports_32; // @[PEArray.scala 74:42]
  assign global_row_pes_0_0_io_in_kv = local_pes_31_0_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_0_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_0_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_0_io_in_stage = io_stage_ports_32; // @[PEArray.scala 75:46]
  assign global_row_pes_0_1_clock = clock;
  assign global_row_pes_0_1_reset = reset;
  assign global_row_pes_0_1_io_in_q = global_row_pes_0_0_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_1_io_in_sum = global_row_pes_0_0_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_1_io_in_sum_exp = 5'sh0; // @[PEArray.scala 77:48]
  assign global_row_pes_0_1_io_in_kv = local_pes_31_1_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_1_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_1_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_1_io_in_stage = global_row_pes_0_0_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_2_clock = clock;
  assign global_row_pes_0_2_reset = reset;
  assign global_row_pes_0_2_io_in_q = global_row_pes_0_1_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_2_io_in_sum = global_row_pes_0_1_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_2_io_in_sum_exp = global_row_pes_0_1_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_2_io_in_kv = local_pes_31_2_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_2_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_2_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_2_io_in_stage = global_row_pes_0_1_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_3_clock = clock;
  assign global_row_pes_0_3_reset = reset;
  assign global_row_pes_0_3_io_in_q = global_row_pes_0_2_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_3_io_in_sum = global_row_pes_0_2_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_3_io_in_sum_exp = global_row_pes_0_2_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_3_io_in_kv = local_pes_31_3_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_3_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_3_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_3_io_in_stage = global_row_pes_0_2_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_4_clock = clock;
  assign global_row_pes_0_4_reset = reset;
  assign global_row_pes_0_4_io_in_q = global_row_pes_0_3_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_4_io_in_sum = global_row_pes_0_3_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_4_io_in_sum_exp = global_row_pes_0_3_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_4_io_in_kv = local_pes_31_4_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_4_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_4_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_4_io_in_stage = global_row_pes_0_3_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_5_clock = clock;
  assign global_row_pes_0_5_reset = reset;
  assign global_row_pes_0_5_io_in_q = global_row_pes_0_4_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_5_io_in_sum = global_row_pes_0_4_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_5_io_in_sum_exp = global_row_pes_0_4_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_5_io_in_kv = local_pes_31_5_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_5_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_5_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_5_io_in_stage = global_row_pes_0_4_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_6_clock = clock;
  assign global_row_pes_0_6_reset = reset;
  assign global_row_pes_0_6_io_in_q = global_row_pes_0_5_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_6_io_in_sum = global_row_pes_0_5_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_6_io_in_sum_exp = global_row_pes_0_5_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_6_io_in_kv = local_pes_31_6_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_6_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_6_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_6_io_in_stage = global_row_pes_0_5_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_7_clock = clock;
  assign global_row_pes_0_7_reset = reset;
  assign global_row_pes_0_7_io_in_q = global_row_pes_0_6_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_7_io_in_sum = global_row_pes_0_6_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_7_io_in_sum_exp = global_row_pes_0_6_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_7_io_in_kv = local_pes_31_7_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_7_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_7_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_7_io_in_stage = global_row_pes_0_6_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_8_clock = clock;
  assign global_row_pes_0_8_reset = reset;
  assign global_row_pes_0_8_io_in_q = global_row_pes_0_7_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_8_io_in_sum = global_row_pes_0_7_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_8_io_in_sum_exp = global_row_pes_0_7_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_8_io_in_kv = local_pes_31_8_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_8_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_8_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_8_io_in_stage = global_row_pes_0_7_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_9_clock = clock;
  assign global_row_pes_0_9_reset = reset;
  assign global_row_pes_0_9_io_in_q = global_row_pes_0_8_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_9_io_in_sum = global_row_pes_0_8_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_9_io_in_sum_exp = global_row_pes_0_8_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_9_io_in_kv = local_pes_31_9_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_9_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_9_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_9_io_in_stage = global_row_pes_0_8_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_10_clock = clock;
  assign global_row_pes_0_10_reset = reset;
  assign global_row_pes_0_10_io_in_q = global_row_pes_0_9_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_10_io_in_sum = global_row_pes_0_9_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_10_io_in_sum_exp = global_row_pes_0_9_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_10_io_in_kv = local_pes_31_10_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_10_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_10_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_10_io_in_stage = global_row_pes_0_9_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_11_clock = clock;
  assign global_row_pes_0_11_reset = reset;
  assign global_row_pes_0_11_io_in_q = global_row_pes_0_10_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_11_io_in_sum = global_row_pes_0_10_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_11_io_in_sum_exp = global_row_pes_0_10_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_11_io_in_kv = local_pes_31_11_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_11_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_11_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_11_io_in_stage = global_row_pes_0_10_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_12_clock = clock;
  assign global_row_pes_0_12_reset = reset;
  assign global_row_pes_0_12_io_in_q = global_row_pes_0_11_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_12_io_in_sum = global_row_pes_0_11_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_12_io_in_sum_exp = global_row_pes_0_11_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_12_io_in_kv = local_pes_31_12_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_12_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_12_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_12_io_in_stage = global_row_pes_0_11_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_13_clock = clock;
  assign global_row_pes_0_13_reset = reset;
  assign global_row_pes_0_13_io_in_q = global_row_pes_0_12_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_13_io_in_sum = global_row_pes_0_12_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_13_io_in_sum_exp = global_row_pes_0_12_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_13_io_in_kv = local_pes_31_13_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_13_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_13_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_13_io_in_stage = global_row_pes_0_12_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_14_clock = clock;
  assign global_row_pes_0_14_reset = reset;
  assign global_row_pes_0_14_io_in_q = global_row_pes_0_13_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_14_io_in_sum = global_row_pes_0_13_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_14_io_in_sum_exp = global_row_pes_0_13_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_14_io_in_kv = local_pes_31_14_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_14_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_14_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_14_io_in_stage = global_row_pes_0_13_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_15_clock = clock;
  assign global_row_pes_0_15_reset = reset;
  assign global_row_pes_0_15_io_in_q = global_row_pes_0_14_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_15_io_in_sum = global_row_pes_0_14_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_15_io_in_sum_exp = global_row_pes_0_14_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_15_io_in_kv = local_pes_31_15_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_15_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_15_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_15_io_in_stage = global_row_pes_0_14_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_16_clock = clock;
  assign global_row_pes_0_16_reset = reset;
  assign global_row_pes_0_16_io_in_q = global_row_pes_0_15_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_16_io_in_sum = global_row_pes_0_15_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_16_io_in_sum_exp = global_row_pes_0_15_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_16_io_in_kv = local_pes_31_16_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_16_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_16_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_16_io_in_stage = global_row_pes_0_15_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_17_clock = clock;
  assign global_row_pes_0_17_reset = reset;
  assign global_row_pes_0_17_io_in_q = global_row_pes_0_16_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_17_io_in_sum = global_row_pes_0_16_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_17_io_in_sum_exp = global_row_pes_0_16_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_17_io_in_kv = local_pes_31_17_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_17_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_17_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_17_io_in_stage = global_row_pes_0_16_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_18_clock = clock;
  assign global_row_pes_0_18_reset = reset;
  assign global_row_pes_0_18_io_in_q = global_row_pes_0_17_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_18_io_in_sum = global_row_pes_0_17_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_18_io_in_sum_exp = global_row_pes_0_17_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_18_io_in_kv = local_pes_31_18_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_18_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_18_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_18_io_in_stage = global_row_pes_0_17_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_19_clock = clock;
  assign global_row_pes_0_19_reset = reset;
  assign global_row_pes_0_19_io_in_q = global_row_pes_0_18_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_19_io_in_sum = global_row_pes_0_18_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_19_io_in_sum_exp = global_row_pes_0_18_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_19_io_in_kv = local_pes_31_19_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_19_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_19_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_19_io_in_stage = global_row_pes_0_18_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_20_clock = clock;
  assign global_row_pes_0_20_reset = reset;
  assign global_row_pes_0_20_io_in_q = global_row_pes_0_19_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_20_io_in_sum = global_row_pes_0_19_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_20_io_in_sum_exp = global_row_pes_0_19_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_20_io_in_kv = local_pes_31_20_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_20_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_20_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_20_io_in_stage = global_row_pes_0_19_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_21_clock = clock;
  assign global_row_pes_0_21_reset = reset;
  assign global_row_pes_0_21_io_in_q = global_row_pes_0_20_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_21_io_in_sum = global_row_pes_0_20_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_21_io_in_sum_exp = global_row_pes_0_20_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_21_io_in_kv = local_pes_31_21_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_21_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_21_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_21_io_in_stage = global_row_pes_0_20_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_22_clock = clock;
  assign global_row_pes_0_22_reset = reset;
  assign global_row_pes_0_22_io_in_q = global_row_pes_0_21_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_22_io_in_sum = global_row_pes_0_21_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_22_io_in_sum_exp = global_row_pes_0_21_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_22_io_in_kv = local_pes_31_22_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_22_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_22_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_22_io_in_stage = global_row_pes_0_21_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_23_clock = clock;
  assign global_row_pes_0_23_reset = reset;
  assign global_row_pes_0_23_io_in_q = global_row_pes_0_22_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_23_io_in_sum = global_row_pes_0_22_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_23_io_in_sum_exp = global_row_pes_0_22_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_23_io_in_kv = local_pes_31_23_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_23_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_23_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_23_io_in_stage = global_row_pes_0_22_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_24_clock = clock;
  assign global_row_pes_0_24_reset = reset;
  assign global_row_pes_0_24_io_in_q = global_row_pes_0_23_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_24_io_in_sum = global_row_pes_0_23_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_24_io_in_sum_exp = global_row_pes_0_23_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_24_io_in_kv = local_pes_31_24_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_24_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_24_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_24_io_in_stage = global_row_pes_0_23_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_25_clock = clock;
  assign global_row_pes_0_25_reset = reset;
  assign global_row_pes_0_25_io_in_q = global_row_pes_0_24_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_25_io_in_sum = global_row_pes_0_24_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_25_io_in_sum_exp = global_row_pes_0_24_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_25_io_in_kv = local_pes_31_25_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_25_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_25_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_25_io_in_stage = global_row_pes_0_24_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_26_clock = clock;
  assign global_row_pes_0_26_reset = reset;
  assign global_row_pes_0_26_io_in_q = global_row_pes_0_25_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_26_io_in_sum = global_row_pes_0_25_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_26_io_in_sum_exp = global_row_pes_0_25_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_26_io_in_kv = local_pes_31_26_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_26_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_26_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_26_io_in_stage = global_row_pes_0_25_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_27_clock = clock;
  assign global_row_pes_0_27_reset = reset;
  assign global_row_pes_0_27_io_in_q = global_row_pes_0_26_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_27_io_in_sum = global_row_pes_0_26_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_27_io_in_sum_exp = global_row_pes_0_26_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_27_io_in_kv = local_pes_31_27_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_27_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_27_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_27_io_in_stage = global_row_pes_0_26_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_28_clock = clock;
  assign global_row_pes_0_28_reset = reset;
  assign global_row_pes_0_28_io_in_q = global_row_pes_0_27_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_28_io_in_sum = global_row_pes_0_27_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_28_io_in_sum_exp = global_row_pes_0_27_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_28_io_in_kv = local_pes_31_28_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_28_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_28_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_28_io_in_stage = global_row_pes_0_27_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_29_clock = clock;
  assign global_row_pes_0_29_reset = reset;
  assign global_row_pes_0_29_io_in_q = global_row_pes_0_28_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_29_io_in_sum = global_row_pes_0_28_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_29_io_in_sum_exp = global_row_pes_0_28_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_29_io_in_kv = local_pes_31_29_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_29_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_29_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_29_io_in_stage = global_row_pes_0_28_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_30_clock = clock;
  assign global_row_pes_0_30_reset = reset;
  assign global_row_pes_0_30_io_in_q = global_row_pes_0_29_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_30_io_in_sum = global_row_pes_0_29_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_30_io_in_sum_exp = global_row_pes_0_29_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_30_io_in_kv = local_pes_31_30_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_30_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_30_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_30_io_in_stage = global_row_pes_0_29_io_out_stage; // @[PEArray.scala 75:46]
  assign global_row_pes_0_31_clock = clock;
  assign global_row_pes_0_31_reset = reset;
  assign global_row_pes_0_31_io_in_q = global_row_pes_0_30_io_out_q; // @[PEArray.scala 74:42]
  assign global_row_pes_0_31_io_in_sum = global_row_pes_0_30_io_out_sum; // @[PEArray.scala 76:44]
  assign global_row_pes_0_31_io_in_sum_exp = global_row_pes_0_30_io_out_sum_exp; // @[PEArray.scala 77:48]
  assign global_row_pes_0_31_io_in_kv = local_pes_31_31_io_out_kv; // @[PEArray.scala 78:43]
  assign global_row_pes_0_31_io_in_inv_sum_exp = inv_modules_32_io_out_inv_sum_exp; // @[PEArray.scala 80:52]
  assign global_row_pes_0_31_io_in_inv_sum = _GEN_2112[8:0]; // @[PEArray.scala 79:48]
  assign global_row_pes_0_31_io_in_stage = global_row_pes_0_30_io_out_stage; // @[PEArray.scala 75:46]
  assign inv_modules_0_io_in_sum = global_col_pes_0_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_0_io_in_exp = global_col_pes_0_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_1_io_in_sum = global_col_pes_1_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_1_io_in_exp = global_col_pes_1_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_2_io_in_sum = global_col_pes_2_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_2_io_in_exp = global_col_pes_2_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_3_io_in_sum = global_col_pes_3_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_3_io_in_exp = global_col_pes_3_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_4_io_in_sum = global_col_pes_4_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_4_io_in_exp = global_col_pes_4_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_5_io_in_sum = global_col_pes_5_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_5_io_in_exp = global_col_pes_5_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_6_io_in_sum = global_col_pes_6_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_6_io_in_exp = global_col_pes_6_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_7_io_in_sum = global_col_pes_7_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_7_io_in_exp = global_col_pes_7_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_8_io_in_sum = global_col_pes_8_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_8_io_in_exp = global_col_pes_8_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_9_io_in_sum = global_col_pes_9_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_9_io_in_exp = global_col_pes_9_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_10_io_in_sum = global_col_pes_10_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_10_io_in_exp = global_col_pes_10_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_11_io_in_sum = global_col_pes_11_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_11_io_in_exp = global_col_pes_11_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_12_io_in_sum = global_col_pes_12_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_12_io_in_exp = global_col_pes_12_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_13_io_in_sum = global_col_pes_13_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_13_io_in_exp = global_col_pes_13_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_14_io_in_sum = global_col_pes_14_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_14_io_in_exp = global_col_pes_14_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_15_io_in_sum = global_col_pes_15_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_15_io_in_exp = global_col_pes_15_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_16_io_in_sum = global_col_pes_16_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_16_io_in_exp = global_col_pes_16_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_17_io_in_sum = global_col_pes_17_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_17_io_in_exp = global_col_pes_17_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_18_io_in_sum = global_col_pes_18_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_18_io_in_exp = global_col_pes_18_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_19_io_in_sum = global_col_pes_19_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_19_io_in_exp = global_col_pes_19_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_20_io_in_sum = global_col_pes_20_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_20_io_in_exp = global_col_pes_20_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_21_io_in_sum = global_col_pes_21_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_21_io_in_exp = global_col_pes_21_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_22_io_in_sum = global_col_pes_22_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_22_io_in_exp = global_col_pes_22_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_23_io_in_sum = global_col_pes_23_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_23_io_in_exp = global_col_pes_23_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_24_io_in_sum = global_col_pes_24_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_24_io_in_exp = global_col_pes_24_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_25_io_in_sum = global_col_pes_25_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_25_io_in_exp = global_col_pes_25_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_26_io_in_sum = global_col_pes_26_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_26_io_in_exp = global_col_pes_26_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_27_io_in_sum = global_col_pes_27_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_27_io_in_exp = global_col_pes_27_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_28_io_in_sum = global_col_pes_28_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_28_io_in_exp = global_col_pes_28_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_29_io_in_sum = global_col_pes_29_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_29_io_in_exp = global_col_pes_29_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_30_io_in_sum = global_col_pes_30_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_30_io_in_exp = global_col_pes_30_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_31_io_in_sum = global_col_pes_31_0_io_out_sum; // @[PEArray.scala 85:34]
  assign inv_modules_31_io_in_exp = global_col_pes_31_0_io_out_sum_exp; // @[PEArray.scala 86:34]
  assign inv_modules_32_io_in_sum = global_row_pes_0_31_io_out_sum; // @[PEArray.scala 90:43]
  assign inv_modules_32_io_in_exp = global_row_pes_0_31_io_out_sum_exp; // @[PEArray.scala 91:43]
  assign weighted_sum_modules_0_clock = clock;
  assign weighted_sum_modules_0_reset = reset;
  assign weighted_sum_modules_0_io_in_sum = global_col_pes_0_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_0_io_in_exp = global_col_pes_0_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_0_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_1_clock = clock;
  assign weighted_sum_modules_1_reset = reset;
  assign weighted_sum_modules_1_io_in_sum = global_col_pes_1_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_1_io_in_exp = global_col_pes_1_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_1_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_2_clock = clock;
  assign weighted_sum_modules_2_reset = reset;
  assign weighted_sum_modules_2_io_in_sum = global_col_pes_2_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_2_io_in_exp = global_col_pes_2_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_2_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_3_clock = clock;
  assign weighted_sum_modules_3_reset = reset;
  assign weighted_sum_modules_3_io_in_sum = global_col_pes_3_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_3_io_in_exp = global_col_pes_3_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_3_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_4_clock = clock;
  assign weighted_sum_modules_4_reset = reset;
  assign weighted_sum_modules_4_io_in_sum = global_col_pes_4_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_4_io_in_exp = global_col_pes_4_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_4_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_5_clock = clock;
  assign weighted_sum_modules_5_reset = reset;
  assign weighted_sum_modules_5_io_in_sum = global_col_pes_5_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_5_io_in_exp = global_col_pes_5_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_5_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_6_clock = clock;
  assign weighted_sum_modules_6_reset = reset;
  assign weighted_sum_modules_6_io_in_sum = global_col_pes_6_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_6_io_in_exp = global_col_pes_6_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_6_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_7_clock = clock;
  assign weighted_sum_modules_7_reset = reset;
  assign weighted_sum_modules_7_io_in_sum = global_col_pes_7_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_7_io_in_exp = global_col_pes_7_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_7_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_8_clock = clock;
  assign weighted_sum_modules_8_reset = reset;
  assign weighted_sum_modules_8_io_in_sum = global_col_pes_8_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_8_io_in_exp = global_col_pes_8_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_8_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_9_clock = clock;
  assign weighted_sum_modules_9_reset = reset;
  assign weighted_sum_modules_9_io_in_sum = global_col_pes_9_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_9_io_in_exp = global_col_pes_9_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_9_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_10_clock = clock;
  assign weighted_sum_modules_10_reset = reset;
  assign weighted_sum_modules_10_io_in_sum = global_col_pes_10_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_10_io_in_exp = global_col_pes_10_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_10_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_11_clock = clock;
  assign weighted_sum_modules_11_reset = reset;
  assign weighted_sum_modules_11_io_in_sum = global_col_pes_11_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_11_io_in_exp = global_col_pes_11_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_11_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_12_clock = clock;
  assign weighted_sum_modules_12_reset = reset;
  assign weighted_sum_modules_12_io_in_sum = global_col_pes_12_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_12_io_in_exp = global_col_pes_12_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_12_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_13_clock = clock;
  assign weighted_sum_modules_13_reset = reset;
  assign weighted_sum_modules_13_io_in_sum = global_col_pes_13_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_13_io_in_exp = global_col_pes_13_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_13_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_14_clock = clock;
  assign weighted_sum_modules_14_reset = reset;
  assign weighted_sum_modules_14_io_in_sum = global_col_pes_14_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_14_io_in_exp = global_col_pes_14_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_14_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_15_clock = clock;
  assign weighted_sum_modules_15_reset = reset;
  assign weighted_sum_modules_15_io_in_sum = global_col_pes_15_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_15_io_in_exp = global_col_pes_15_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_15_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_16_clock = clock;
  assign weighted_sum_modules_16_reset = reset;
  assign weighted_sum_modules_16_io_in_sum = global_col_pes_16_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_16_io_in_exp = global_col_pes_16_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_16_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_17_clock = clock;
  assign weighted_sum_modules_17_reset = reset;
  assign weighted_sum_modules_17_io_in_sum = global_col_pes_17_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_17_io_in_exp = global_col_pes_17_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_17_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_18_clock = clock;
  assign weighted_sum_modules_18_reset = reset;
  assign weighted_sum_modules_18_io_in_sum = global_col_pes_18_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_18_io_in_exp = global_col_pes_18_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_18_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_19_clock = clock;
  assign weighted_sum_modules_19_reset = reset;
  assign weighted_sum_modules_19_io_in_sum = global_col_pes_19_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_19_io_in_exp = global_col_pes_19_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_19_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_20_clock = clock;
  assign weighted_sum_modules_20_reset = reset;
  assign weighted_sum_modules_20_io_in_sum = global_col_pes_20_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_20_io_in_exp = global_col_pes_20_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_20_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_21_clock = clock;
  assign weighted_sum_modules_21_reset = reset;
  assign weighted_sum_modules_21_io_in_sum = global_col_pes_21_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_21_io_in_exp = global_col_pes_21_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_21_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_22_clock = clock;
  assign weighted_sum_modules_22_reset = reset;
  assign weighted_sum_modules_22_io_in_sum = global_col_pes_22_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_22_io_in_exp = global_col_pes_22_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_22_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_23_clock = clock;
  assign weighted_sum_modules_23_reset = reset;
  assign weighted_sum_modules_23_io_in_sum = global_col_pes_23_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_23_io_in_exp = global_col_pes_23_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_23_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_24_clock = clock;
  assign weighted_sum_modules_24_reset = reset;
  assign weighted_sum_modules_24_io_in_sum = global_col_pes_24_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_24_io_in_exp = global_col_pes_24_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_24_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_25_clock = clock;
  assign weighted_sum_modules_25_reset = reset;
  assign weighted_sum_modules_25_io_in_sum = global_col_pes_25_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_25_io_in_exp = global_col_pes_25_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_25_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_26_clock = clock;
  assign weighted_sum_modules_26_reset = reset;
  assign weighted_sum_modules_26_io_in_sum = global_col_pes_26_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_26_io_in_exp = global_col_pes_26_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_26_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_27_clock = clock;
  assign weighted_sum_modules_27_reset = reset;
  assign weighted_sum_modules_27_io_in_sum = global_col_pes_27_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_27_io_in_exp = global_col_pes_27_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_27_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_28_clock = clock;
  assign weighted_sum_modules_28_reset = reset;
  assign weighted_sum_modules_28_io_in_sum = global_col_pes_28_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_28_io_in_exp = global_col_pes_28_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_28_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_29_clock = clock;
  assign weighted_sum_modules_29_reset = reset;
  assign weighted_sum_modules_29_io_in_sum = global_col_pes_29_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_29_io_in_exp = global_col_pes_29_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_29_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_30_clock = clock;
  assign weighted_sum_modules_30_reset = reset;
  assign weighted_sum_modules_30_io_in_sum = global_col_pes_30_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_30_io_in_exp = global_col_pes_30_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_30_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_31_clock = clock;
  assign weighted_sum_modules_31_reset = reset;
  assign weighted_sum_modules_31_io_in_sum = global_col_pes_31_0_io_out_sum; // @[PEArray.scala 95:43]
  assign weighted_sum_modules_31_io_in_exp = global_col_pes_31_0_io_out_sum_exp; // @[PEArray.scala 96:43]
  assign weighted_sum_modules_31_io_control = io_weight_control; // @[PEArray.scala 97:44]
  assign weighted_sum_modules_32_clock = clock;
  assign weighted_sum_modules_32_reset = reset;
  assign weighted_sum_modules_32_io_in_sum = global_row_pes_0_31_io_out_sum; // @[PEArray.scala 102:52]
  assign weighted_sum_modules_32_io_in_exp = global_row_pes_0_31_io_out_sum_exp; // @[PEArray.scala 103:52]
  assign weighted_sum_modules_32_io_control = io_weight_control; // @[PEArray.scala 104:53]
endmodule
